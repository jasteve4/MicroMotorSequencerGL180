* NGSPICE file created from driver_core.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

.subckt driver_core clock clock_a col_select_a[0] col_select_a[1] col_select_a[2]
+ col_select_a[3] col_select_a[4] col_select_a[5] data_in_a[0] data_in_a[10] data_in_a[11]
+ data_in_a[12] data_in_a[13] data_in_a[14] data_in_a[15] data_in_a[1] data_in_a[2]
+ data_in_a[3] data_in_a[4] data_in_a[5] data_in_a[6] data_in_a[7] data_in_a[8] data_in_a[9]
+ driver_io[0] driver_io[1] inverter_select_a mem_address_a[0] mem_address_a[1] mem_address_a[2]
+ mem_address_a[3] mem_address_a[4] mem_address_a[5] mem_address_a[6] mem_address_a[7]
+ mem_address_a[8] mem_address_a[9] mem_write_n_a output_active_a row_col_select_a
+ row_select_a[0] row_select_a[1] row_select_a[2] row_select_a[3] row_select_a[4]
+ row_select_a[5] vccd1 vssd1
XFILLER_39_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07383__I _02611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11705__I1 u2.mem\[181\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06883_ _02338_ _02345_ _02362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09671_ _04550_ _00582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06337__A2 _01834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12595__CLK clknet_leaf_105_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07534__A1 _03002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08622_ _03808_ u2.mem\[12\]\[4\] _03885_ _03886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06888__A3 _02344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08553_ _03845_ _00169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07504_ u2.mem\[1\]\[7\] _02795_ _02796_ u2.mem\[7\]\[7\] _02976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07298__B1 _02688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08484_ _03799_ _03800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_35_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07435_ u2.mem\[29\]\[5\] _02833_ _02834_ u2.mem\[11\]\[5\] _02909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10841__A1 _03983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07366_ u2.mem\[28\]\[4\] _02839_ _02840_ u2.mem\[31\]\[4\] _02841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08637__I1 u2.mem\[12\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_350_clock clknet_5_4_0_clock clknet_leaf_350_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_143_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09105_ _04199_ _00367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06317_ u2.mem\[158\]\[3\] _01728_ _01729_ u2.mem\[151\]\[3\] _01731_ u2.mem\[193\]\[3\]
+ _01821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_52_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07297_ _02769_ _02770_ _02771_ _02772_ _02773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_163_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07558__I _02470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09036_ _04152_ _00345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07470__B1 _02888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06248_ _01597_ _01754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06462__I _01914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06179_ _01563_ _01677_ _01587_ _01686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_172_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06025__A1 _01516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13370__CLK clknet_leaf_357_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06576__A2 _02053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10712__I _05195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09938_ _04689_ u2.mem\[42\]\[3\] _04719_ _04723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07507__B _02978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09869_ _04605_ u2.mem\[40\]\[12\] _04676_ _04677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06328__A2 _01712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07525__B2 u2.mem\[10\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11900_ _05927_ _05942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_133_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12880_ _00759_ clknet_leaf_230_clock u2.mem\[47\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_303_clock clknet_5_16_0_clock clknet_leaf_303_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11831_ _05870_ u2.mem\[189\]\[2\] _05896_ _05899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07540__A4 _03011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07289__B1 _02570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11762_ _04248_ _05847_ _05856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_60_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09013__I data_in_trans\[3\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13501_ _01380_ clknet_leaf_330_clock u2.mem\[187\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10713_ _05194_ u2.mem\[61\]\[0\] _05196_ _05197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12318__CLK clknet_leaf_199_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11880__I0 u2.mem\[192\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11693_ _05794_ u2.mem\[180\]\[3\] _05810_ _05814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13432_ _01311_ clknet_leaf_336_clock u2.mem\[175\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_318_clock clknet_5_18_0_clock clknet_leaf_318_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08852__I _03692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10644_ _05156_ _00949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08628__I1 u2.mem\[12\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11632__I0 _05756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10575_ _05114_ _00922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13363_ _01242_ clknet_leaf_358_clock u2.mem\[164\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12314_ _00193_ clknet_leaf_118_clock u2.mem\[11\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12468__CLK clknet_leaf_105_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13294_ _01173_ clknet_leaf_364_clock u2.mem\[152\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12026__D row_select_trans\[0\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11919__S _05950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08005__A2 _03464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12245_ _00124_ clknet_leaf_73_clock u2.mem\[7\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07213__B1 _02614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11935__I1 u2.mem\[193\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12176_ _00055_ clknet_leaf_226_clock u2.mem\[3\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11718__I _03662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07764__B2 u2.mem\[25\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11127_ _05457_ _01131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08299__I _03674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11058_ _05384_ u2.mem\[141\]\[1\] _05413_ _05415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08564__I0 _03826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07516__B2 u2.mem\[46\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10009_ _04685_ u2.mem\[44\]\[1\] _04762_ _04764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_76_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07819__A2 _03269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11871__I0 _05915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06991__B _02468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13243__CLK clknet_leaf_291_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07220_ u2.mem\[40\]\[2\] _02406_ _02415_ u2.mem\[30\]\[2\] _02697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08619__I1 u2.mem\[12\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07151_ u2.mem\[5\]\[0\] _02627_ _02629_ u2.mem\[38\]\[0\] _02630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_67_clock_I clknet_5_9_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09292__I1 u2.mem\[27\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06102_ _01547_ _01608_ _01609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_146_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09794__S _04633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06255__B2 u2.mem\[153\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07082_ _02560_ _02561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13393__CLK clknet_5_16_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11829__S _05896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06033_ _01528_ _01540_ _01541_ _01542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07204__B1 _02681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11926__I1 u2.mem\[193\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07327__B _02745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07984_ u2.mem\[17\]\[15\] _03310_ _03311_ u2.mem\[24\]\[15\] _03448_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09723_ data_in_trans\[6\].data_sync _04585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06935_ _02407_ _02408_ _02411_ _02413_ _02414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__07046__C _02394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08555__I0 _03817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11564__S _05731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09654_ _04496_ u2.mem\[35\]\[14\] _04537_ _04540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06866_ _02339_ _02344_ _02345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08605_ _03831_ u2.mem\[11\]\[14\] _03872_ _03875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09585_ _04500_ _04501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06797_ u2.mem\[164\]\[4\] _02050_ _02054_ u2.mem\[178\]\[4\] _02278_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08307__I0 _03681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09969__S _04740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08536_ _03835_ _03836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08873__S _04042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_344_clock_I clknet_5_5_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08467_ _03698_ u2.mem\[8\]\[9\] _03788_ _03790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10908__S _05319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08483__A2 _03544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07418_ u2.mem\[14\]\[5\] _02890_ _02891_ u2.mem\[12\]\[5\] _02892_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08398_ _03723_ u2.mem\[6\]\[15\] _03743_ _03747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12610__CLK clknet_leaf_173_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11614__I0 _05754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07349_ u2.mem\[60\]\[4\] _02822_ _02823_ u2.mem\[62\]\[4\] _02824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06246__A1 u2.mem\[159\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10360_ _04978_ _00843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06192__I _01698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06246__B2 u2.mem\[149\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07994__A1 _01980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11739__S _05840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09019_ _04138_ _04139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10291_ _04913_ u2.mem\[50\]\[12\] _04938_ _04939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10643__S _05152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06261__A4 _01766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12030_ row_select_trans\[2\].A clknet_leaf_307_clock row_select_trans\[2\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11917__I1 u2.mem\[193\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09209__S _04261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06920__I _02370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06549__A2 _02033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09008__I data_in_trans\[2\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13116__CLK clknet_leaf_261_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08546__I0 _03808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12932_ _00811_ clknet_leaf_66_clock u2.mem\[50\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_242_clock clknet_5_19_0_clock clknet_leaf_242_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12863_ _00742_ clknet_leaf_148_clock u2.mem\[46\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12140__CLK clknet_leaf_211_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06721__A2 _01995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13266__CLK clknet_leaf_295_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11814_ _05889_ _01386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12794_ _00673_ clknet_leaf_48_clock u2.mem\[41\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_257_clock clknet_5_23_0_clock clknet_leaf_257_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11745_ _05837_ u2.mem\[183\]\[5\] _05839_ _05846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09678__I _04543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08582__I _03856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07700__B _02978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12290__CLK clknet_leaf_165_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11676_ _05792_ u2.mem\[179\]\[2\] _05801_ _05804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13415_ _01294_ clknet_leaf_342_clock u2.mem\[172\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10627_ _05121_ u2.mem\[58\]\[12\] _05146_ _05147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10617__I _05130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07434__B1 _02907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13346_ _01225_ clknet_leaf_5_clock u2.mem\[161\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10558_ _05102_ _00917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06788__A2 _02267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13277_ _01156_ clknet_leaf_10_clock u2.mem\[149\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10489_ _05050_ _05061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_29_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12228_ _00107_ clknet_leaf_64_clock u2.mem\[6\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07737__A1 u2.mem\[40\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07737__B2 u2.mem\[30\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07147__B _02484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12159_ _00038_ clknet_leaf_153_clock u2.mem\[2\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08958__S _04097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_293_clock_I clknet_5_20_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08537__I0 _03798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06720_ _02179_ _02190_ _02194_ _02203_ _02204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_65_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06651_ _02119_ _02044_ _02136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09789__S _04628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09370_ _04363_ _00468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06582_ _02045_ _02018_ _02067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12633__CLK clknet_leaf_103_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08321_ _03692_ _03693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08252_ _03642_ _00071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07673__B1 _03070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07203_ _02597_ _02681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08183_ _03599_ _00045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10527__I _05072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12783__CLK clknet_leaf_322_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07134_ _02466_ _02467_ _02498_ _02394_ _02613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_88_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11221__A1 _05354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06779__A2 _02042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07065_ _02347_ _02544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07836__I _02581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12013__CLK clknet_2_0__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06016_ u2.driver_mem\[5\] _01518_ _01525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__13139__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07728__B2 u2.mem\[38\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11524__A2 _05690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10583__I0 _05119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input36_I row_col_select_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06400__A1 u2.mem\[144\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06400__B2 u2.mem\[182\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07967_ u2.mem\[44\]\[15\] _02521_ _02523_ u2.mem\[42\]\[15\] _03431_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12163__CLK clknet_leaf_91_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11294__S _05558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09706_ _04130_ _04572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06918_ u2.mem\[32\]\[0\] _02386_ _02396_ u2.mem\[2\]\[0\] _02397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08667__I _03905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07898_ u2.mem\[17\]\[13\] _03310_ _03311_ u2.mem\[24\]\[13\] _03364_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07571__I _02494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09637_ _04530_ _00568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06849_ u2.mem\[154\]\[5\] _02225_ _02226_ u2.mem\[162\]\[5\] _02328_ _02329_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_55_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06187__I _01693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09568_ _04163_ _04489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08519_ _03705_ _03824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11835__I0 _05874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09499_ _04445_ _00515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07259__A3 _02730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08700__I0 _03937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11530_ _05712_ _01279_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07664__B1 _03133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06915__I _02363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11461_ _05667_ _05668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13200_ _01079_ clknet_leaf_271_clock u2.mem\[136\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06219__A1 _01545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10412_ _05014_ u2.mem\[53\]\[9\] _05012_ _05015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11392_ _05295_ _05606_ _05624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_152_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13131_ _01010_ clknet_leaf_246_clock u2.mem\[63\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10343_ _04891_ u2.mem\[52\]\[2\] _04966_ _04969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10274_ _04929_ _00806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13062_ _00941_ clknet_leaf_30_clock u2.mem\[58\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07982__A4 _03445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07719__A1 u2.mem\[29\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12506__CLK clknet_leaf_121_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12013_ net28 clknet_2_0__leaf_clock_a mem_address_trans\[4\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10574__I0 _05112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_181_clock clknet_5_30_0_clock clknet_leaf_181_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_15_clock_I clknet_5_2_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12656__CLK clknet_leaf_221_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12915_ _00794_ clknet_leaf_147_clock u2.mem\[49\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06155__C2 u2.mem\[181\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06097__I _01603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_196_clock clknet_5_31_0_clock clknet_leaf_196_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12846_ _00725_ clknet_leaf_203_clock u2.mem\[45\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12777_ _00656_ clknet_leaf_130_clock u2.mem\[40\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10548__S _05095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07655__B1 _03124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11728_ _05835_ u2.mem\[182\]\[4\] _05826_ _05836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09201__I _04135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10347__I _04965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11659_ _05792_ u2.mem\[178\]\[2\] _05788_ _05793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06046__B _01552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12036__CLK clknet_leaf_311_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11379__S _05616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13329_ _01208_ clknet_leaf_3_clock u2.mem\[158\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_134_clock clknet_5_12_0_clock clknet_leaf_134_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_127_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07656__I _02530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06560__I _02044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12186__CLK clknet_leaf_59_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08870_ _04044_ u2.mem\[17\]\[13\] _04042_ _04045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13431__CLK clknet_leaf_36_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07821_ _02545_ _03288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_149_clock clknet_5_24_0_clock clknet_leaf_149_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_29_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10810__I _05252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08487__I _03663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07752_ u2.mem\[14\]\[11\] _03123_ _03124_ u2.mem\[12\]\[11\] _03220_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06703_ _02101_ _02187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07683_ _02626_ _03153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08930__I0 _04026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11842__S _05905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09422_ _04399_ _00484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06697__A1 u2.mem\[167\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06697__B2 u2.mem\[183\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06634_ _02027_ _02017_ _02119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09353_ _04352_ _00462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11817__I0 _05870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06565_ _02031_ _02041_ _02050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08304_ _03510_ _03679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06449__A1 _01878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06449__B2 _01944_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07646__B1 _03115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09284_ _04311_ _04250_ _04312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_20_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06496_ _01981_ _01927_ _01982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09111__I _04202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08235_ mem_address_trans\[2\].data_sync _03631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07661__A3 _03119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08166_ _03584_ _03590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_162_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12529__CLK clknet_leaf_166_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07117_ _02595_ _02596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08097_ _03479_ _03540_ _03541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_49_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07048_ _02407_ _02408_ _02519_ _02454_ _02527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__06621__A1 u2.mem\[188\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06621__B2 u2.mem\[175\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08598__S _03867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12679__CLK clknet_leaf_130_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08999_ _04121_ _04122_ _04123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_9_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_189_clock_I clknet_5_31_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10961_ _05354_ _05317_ _05355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_56_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11752__S _05849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08921__I0 _04017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12700_ _00579_ clknet_leaf_256_clock u2.mem\[36\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06688__A1 u2.mem\[151\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06688__B2 u2.mem\[158\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10892_ _05309_ _05310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09222__S _04270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12631_ _00510_ clknet_leaf_114_clock u2.mem\[31\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11808__I0 _05876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_241_clock_I clknet_5_19_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07637__B1 _03029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12059__CLK clknet_2_1__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12562_ _00441_ clknet_leaf_171_clock u2.mem\[27\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09021__I _04123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11513_ _05668_ u2.mem\[169\]\[1\] _05700_ _05702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12493_ _00372_ clknet_leaf_186_clock u2.mem\[23\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_51_clock clknet_5_13_0_clock clknet_leaf_51_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11444_ _05627_ u2.mem\[165\]\[1\] _05655_ _05657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11199__S _05502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13454__CLK clknet_leaf_300_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11375_ _05595_ u2.mem\[160\]\[5\] _05607_ _05614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13114_ _00993_ clknet_leaf_333_clock u2.mem\[61\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10326_ _04958_ _00829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_66_clock clknet_5_3_0_clock clknet_leaf_66_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13045_ _00924_ clknet_leaf_25_clock u2.mem\[57\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10257_ _04918_ u2.mem\[49\]\[14\] _04914_ _04919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10188_ _04873_ _00776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10172__A1 _03983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11662__S _05788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06679__A1 _01545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07876__B1 _02505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09132__S _04213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07340__A2 _02660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12829_ _00708_ clknet_leaf_207_clock u2.mem\[44\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11461__I _05667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07891__A3 _03355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06350_ _01849_ _01850_ _01851_ _01852_ _01853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_163_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06281_ u2.mem\[175\]\[2\] _01602_ _01631_ u2.mem\[188\]\[2\] _01786_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06300__B1 _01680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_19_clock clknet_5_2_0_clock clknet_leaf_19_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_102_1511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08020_ mem_address_trans\[1\].data_sync _03481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08770__I _03962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07386__I _02621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06603__A1 _01992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09971_ _04685_ u2.mem\[43\]\[1\] _04740_ _04742_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12821__CLK clknet_leaf_83_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11837__S _05895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08922_ _04076_ _00307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08853_ _04014_ _04033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_131_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08211__S _03614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06367__B1 _01688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06906__A2 _02371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_190_clock_I clknet_5_31_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07804_ u2.mem\[54\]\[12\] _03114_ _03115_ u2.mem\[55\]\[12\] _03271_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_3609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08784_ _03987_ _03988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05996_ u2.select_mem_col\[0\] _01505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07735_ u2.mem\[45\]\[11\] _03099_ _03100_ u2.mem\[34\]\[11\] _03203_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08945__I _04073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07666_ u2.mem\[37\]\[9\] _03058_ _03059_ u2.mem\[59\]\[9\] _03136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12201__CLK clknet_leaf_54_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13327__CLK clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09405_ _04387_ u2.mem\[29\]\[13\] _04385_ _04388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06617_ u2.mem\[187\]\[0\] _02100_ _02101_ u2.mem\[192\]\[0\] _02102_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07597_ u2.mem\[29\]\[8\] _03066_ _03067_ u2.mem\[11\]\[8\] _03068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_94_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09336_ _04263_ u2.mem\[28\]\[5\] _04341_ _04343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07619__B1 _03089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06548_ _02032_ _02011_ _02033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09267_ _04272_ u2.mem\[26\]\[9\] _04300_ _04302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12351__CLK clknet_leaf_148_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10916__S _05318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13477__CLK clknet_leaf_298_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06479_ _01966_ _01955_ _01967_ _01968_ _01460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_166_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08680__I _03905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08218_ _03566_ u2.mem\[3\]\[9\] _03619_ _03621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06842__A1 u2.mem\[145\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06842__B2 u2.mem\[168\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09198_ _04131_ _04256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08149_ _03578_ _00032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10715__I _04991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11160_ _05468_ u2.mem\[147\]\[3\] _05475_ _05479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10111_ _04828_ _00744_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11091_ _05436_ _01116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06070__A2 _01576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09395__I0 _04380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10042_ _04564_ _04782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07570__A2 _03039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06373__A3 _01862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11993_ _00005_ clknet_leaf_318_clock u2.mem\[0\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11482__S _05683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10944_ _04130_ _05342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11281__I _05516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10875_ _05298_ _01038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12614_ _00493_ clknet_leaf_93_clock u2.mem\[30\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08791__S _03990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12545_ _00424_ clknet_leaf_168_clock u2.mem\[26\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12029__D net39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10826__S _05263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06833__A1 u2.mem\[180\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12476_ _00355_ clknet_leaf_181_clock u2.mem\[22\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06833__B2 u2.mem\[172\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11427_ _05646_ _05647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_137_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11358_ _05603_ _01216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10309_ _04943_ _04949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_113_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12994__CLK clknet_leaf_236_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11289_ _05561_ _01189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13028_ _00907_ clknet_leaf_31_clock u2.mem\[56\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11193__I0 _05472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12224__CLK clknet_leaf_231_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07520_ u2.mem\[61\]\[7\] _02899_ _02900_ u2.mem\[63\]\[7\] _02992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_78_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07451_ u2.mem\[6\]\[5\] _02861_ _02862_ u2.mem\[47\]\[5\] _02925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12374__CLK clknet_leaf_78_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07864__A3 _03319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06402_ u2.mem\[170\]\[5\] _01686_ _01688_ u2.mem\[156\]\[5\] _01904_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11248__I1 u2.mem\[152\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07382_ u2.mem\[39\]\[4\] _02855_ _02856_ u2.mem\[48\]\[4\] _02857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09310__I0 _04276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09121_ _04140_ u2.mem\[23\]\[4\] _04208_ _04209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06333_ u2.mem\[191\]\[3\] _01682_ _01684_ u2.mem\[179\]\[3\] _01837_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_137_clock_I clknet_5_13_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06285__C1 u2.mem\[165\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09052_ _04164_ u2.mem\[21\]\[11\] _04155_ _04165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06824__A1 _01844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06264_ _01768_ _01769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_163_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08003_ u2.active_mem\[8\] _03458_ _03459_ u2.active_mem\[9\] _03466_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06195_ _01561_ _01563_ _01580_ _01702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_102_1374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09954_ _04705_ u2.mem\[42\]\[10\] _04729_ _04732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07844__I _02592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08905_ _04065_ _00301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09885_ _04572_ _04687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08836_ _03671_ _04021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08876__S _04042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07552__A2 _03021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08767_ _03976_ _00252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12717__CLK clknet_leaf_254_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07718_ u2.mem\[26\]\[10\] _03139_ _03140_ u2.mem\[10\]\[10\] _03187_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11636__A1 _05285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08698_ _03936_ _00223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07304__A2 _02361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07649_ _03113_ _03116_ _03117_ _03118_ _03119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_53_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06409__B _01910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10660_ _05165_ _00956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12867__CLK clknet_leaf_60_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09301__I0 _04267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09319_ _04285_ u2.mem\[27\]\[15\] _04328_ _04332_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10646__S _05157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10591_ _05125_ _00927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10998__I0 _05346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12330_ _00209_ clknet_leaf_125_clock u2.mem\[12\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06815__A1 u2.mem\[194\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06815__B2 u2.mem\[190\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08116__S _03555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12261_ _00140_ clknet_leaf_70_clock u2.mem\[8\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11212_ _05512_ _01161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12192_ _00071_ clknet_leaf_228_clock u2.mem\[4\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11143_ _05345_ _05468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12247__CLK clknet_leaf_55_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11074_ _05424_ u2.mem\[142\]\[1\] _05422_ _05425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11175__I0 _05468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10025_ _04700_ u2.mem\[44\]\[8\] _04772_ _04773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10922__I0 _05294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07543__A2 _02866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12397__CLK clknet_leaf_180_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06751__B1 _02152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11478__I1 u2.mem\[166\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11976_ _05218_ u2.mem\[194\]\[10\] _05985_ _05986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09540__I0 _04469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10927_ _05330_ _01058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10858_ _05194_ u2.mem\[129\]\[0\] _05287_ _05288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13577_ _01456_ clknet_leaf_35_clock u2.mem\[194\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10789_ _05220_ u2.mem\[62\]\[11\] _05242_ _05246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06806__A1 u2.mem\[180\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12528_ _00407_ clknet_leaf_169_clock u2.mem\[25\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06806__B2 u2.mem\[172\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07074__A4 _02552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12459_ _00338_ clknet_leaf_179_clock u2.mem\[21\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13022__CLK clknet_leaf_259_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11387__S _05615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10291__S _04938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07231__A1 u2.mem\[58\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06034__A2 _01542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07231__B2 u2.mem\[36\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13172__CLK clknet_leaf_263_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06951_ _02369_ _02430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09670_ _04473_ u2.mem\[36\]\[4\] _04549_ _04550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06882_ _02360_ _02361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_63_clock_I clknet_5_9_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08621_ _03879_ _03885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_94_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11914__I _05949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08552_ _03815_ u2.mem\[10\]\[7\] _03841_ _03845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07503_ u2.mem\[15\]\[7\] _02792_ _02793_ u2.mem\[13\]\[7\] _02975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_78_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08483_ _03658_ _03544_ _03776_ _03799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_74_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07434_ u2.mem\[26\]\[5\] _02906_ _02907_ u2.mem\[10\]\[5\] _02908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_165_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07365_ _02586_ _02840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_15_0_clock clknet_3_7_0_clock clknet_4_15_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_clkbuf_leaf_288_clock_I clknet_5_20_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10466__S _05045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07839__I _02586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09104_ _04171_ u2.mem\[22\]\[13\] _04197_ _04199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06258__C1 u2.mem\[172\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06316_ u2.mem\[177\]\[3\] _01734_ _01646_ u2.mem\[165\]\[3\] u2.mem\[163\]\[3\]
+ _01642_ _01820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_143_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06743__I _02127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07296_ u2.mem\[18\]\[3\] _02606_ _02608_ u2.mem\[19\]\[3\] _02772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09035_ _04151_ u2.mem\[21\]\[7\] _04141_ _04152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06247_ _01592_ _01753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07470__B2 u2.mem\[42\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06178_ u2.mem\[191\]\[0\] _01682_ _01684_ u2.mem\[179\]\[0\] _01685_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_132_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_340_clock_I clknet_5_5_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07773__A2 _03088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09937_ _04722_ _00676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09868_ _04660_ _04676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07525__A2 _02906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08819_ _04008_ _00272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09799_ _04636_ _00624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11830_ _05898_ _01393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07289__A1 u2.mem\[29\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11761_ _05855_ _01367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11760__S _05848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13500_ _01379_ clknet_leaf_317_clock u2.mem\[186\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10712_ _05195_ _05196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11692_ _05813_ _01340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11880__I1 _03497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13431_ _01310_ clknet_leaf_36_clock u2.mem\[175\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10643_ _05101_ u2.mem\[59\]\[3\] _05152_ _05156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13045__CLK clknet_leaf_25_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13362_ _01241_ clknet_leaf_354_clock u2.mem\[163\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10574_ _05112_ u2.mem\[57\]\[8\] _05113_ _05114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12313_ _00192_ clknet_leaf_118_clock u2.mem\[11\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13293_ _01172_ clknet_leaf_364_clock u2.mem\[152\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12244_ _00123_ clknet_leaf_74_clock u2.mem\[7\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12175_ _00054_ clknet_leaf_218_clock u2.mem\[3\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07213__B2 u2.mem\[4\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11000__S _05372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07764__A2 _03069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11126_ _05428_ u2.mem\[145\]\[3\] _05453_ _05457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11057_ _05414_ _01104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07516__A2 _02893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08564__I1 u2.mem\[10\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10008_ _04763_ _00706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09204__I _04139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11959_ _05976_ _01444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07819__A3 _03278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11871__I1 u2.mem\[191\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10286__S _04933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07150_ _02628_ _02629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12412__CLK clknet_leaf_198_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13538__CLK clknet_leaf_34_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06101_ _01584_ _01559_ _01608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07081_ _02473_ _02399_ _02400_ _02453_ _02560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_103_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06032_ u2.select_mem_row\[3\] u2.select_mem_col\[3\] _01510_ _01541_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11387__I0 _05593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07983_ u2.mem\[23\]\[15\] _02596_ _02598_ u2.mem\[22\]\[15\] _03447_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11845__S _05905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09722_ _04584_ _00599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06934_ _02412_ _02413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_68_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09653_ _04539_ _00575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06865_ _02340_ _02341_ _02342_ _02343_ _02344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_167_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08604_ _03874_ _00191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09584_ _03583_ _04441_ _04500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_103_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06796_ _02273_ _02274_ _02275_ _02276_ _02277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08535_ _03658_ _03726_ _03776_ _03835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_24_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11311__I0 _05556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13068__CLK clknet_leaf_254_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11580__S _05739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08466_ _03789_ _00138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08483__A3 _03776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07417_ _02527_ _02891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07691__A1 _01958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10196__S _04875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08397_ _03746_ _00112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07569__I _02488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12092__CLK clknet_leaf_302_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06473__I _01913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07348_ _02548_ _02823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08491__I0 _03804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07443__B2 u2.mem\[21\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07279_ u2.mem\[49\]\[3\] _02660_ _02661_ u2.mem\[46\]\[3\] _02755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10924__S _05327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12905__CLK clknet_leaf_141_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09784__I _04617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07994__A2 _03246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09018_ data_in_trans\[4\].data_sync _04138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10290_ _04922_ _04938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_88_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07746__A2 _03111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09991__I0 _04705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08546__I1 u2.mem\[10\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09225__S _04270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12931_ _00810_ clknet_leaf_232_clock u2.mem\[50\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12862_ _00741_ clknet_leaf_199_clock u2.mem\[46\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09024__I data_in_trans\[5\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11813_ _05864_ u2.mem\[188\]\[0\] _05888_ _05889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12793_ _00672_ clknet_leaf_48_clock u2.mem\[41\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11490__S _05682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11744_ _05845_ _01360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12435__CLK clknet_leaf_108_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07682__A1 _03148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11675_ _05803_ _01333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13414_ _01293_ clknet_leaf_342_clock u2.mem\[172\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_11_clock_I clknet_5_3_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10626_ _05130_ _05146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_161_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07029__A4 _02507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07434__A1 u2.mem\[26\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12037__D net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13345_ _01224_ clknet_leaf_4_clock u2.mem\[161\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06237__A2 _01741_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07434__B2 u2.mem\[10\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12585__CLK clknet_leaf_115_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10557_ _05101_ u2.mem\[57\]\[3\] _05095_ _05102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13276_ _01155_ clknet_leaf_11_clock u2.mem\[149\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11369__I0 _05589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10488_ _05060_ _00889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12227_ _00106_ clknet_leaf_64_clock u2.mem\[6\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07198__B1 _02570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09982__I0 _04696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12158_ _00037_ clknet_leaf_205_clock u2.mem\[2\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07147__C _02364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_236_clock_I clknet_5_19_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11665__S _05787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11109_ _05447_ _01123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12089_ net35 clknet_2_0__leaf_clock_a output_active_trans.A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09734__I0 _04592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11464__I _03499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11541__I0 _05719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13210__CLK clknet_leaf_281_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06558__I _02042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06650_ u2.mem\[194\]\[0\] _02133_ _02134_ u2.mem\[190\]\[0\] _02135_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_65_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06581_ _02065_ _02066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_364_clock clknet_5_0_0_clock clknet_leaf_364_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_127_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08320_ _03691_ _03692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13360__CLK clknet_leaf_356_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08251_ _03557_ u2.mem\[4\]\[5\] _03640_ _03642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07673__B2 u2.mem\[25\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12928__CLK clknet_leaf_235_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07202_ _02595_ _02680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08182_ _03570_ u2.mem\[2\]\[11\] _03595_ _03599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07133_ _02611_ _02612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11221__A2 _05482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07064_ u2.mem\[37\]\[0\] _02540_ _02542_ u2.mem\[59\]\[0\] _02543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_145_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_302_clock clknet_5_16_0_clock clknet_leaf_302_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_47_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06015_ u2.driver_mem\[6\] _01513_ _01523_ _01524_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08225__I0 _03572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07728__A2 _03153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09973__I0 _04687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12308__CLK clknet_leaf_100_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06400__A2 _01670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07966_ _03426_ _03427_ _03428_ _03429_ _03430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_114_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_317_clock clknet_5_18_0_clock clknet_leaf_317_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_60_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09705_ _04571_ _00595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09725__I0 _04586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06917_ _02395_ _02396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input29_I mem_address_a[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07897_ u2.mem\[23\]\[13\] _02596_ _02598_ u2.mem\[22\]\[13\] _03363_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11532__I0 _05713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09636_ _04478_ u2.mem\[35\]\[6\] _04527_ _04530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_1568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06848_ _02325_ _02326_ _02327_ _02328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_55_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06468__I _01927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08884__S _04051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12458__CLK clknet_leaf_127_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09567_ _04488_ _00540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06779_ u2.mem\[180\]\[3\] _02042_ _02013_ u2.mem\[172\]\[3\] _02261_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10099__I0 _04786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08518_ _03823_ _00156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08683__I _03697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07801__B _03211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09498_ _04360_ u2.mem\[32\]\[1\] _04443_ _04445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11835__I1 u2.mem\[189\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07259__A4 _02735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08449_ _03664_ u2.mem\[8\]\[1\] _03778_ _03780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10718__I _04994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06467__A2 _01929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11460_ _03496_ _05667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_185_clock_I clknet_5_30_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10411_ _03696_ _05014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11391_ _05499_ _05623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07967__A2 _02521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13130_ _01009_ clknet_leaf_327_clock u2.mem\[62\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10342_ _04968_ _00835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08216__I0 _03563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13061_ _00940_ clknet_leaf_26_clock u2.mem\[58\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10273_ _04895_ u2.mem\[50\]\[4\] _04928_ _04929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07719__A2 _03066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09019__I _04138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12012_ mem_address_trans\[3\].A clknet_leaf_244_clock mem_address_trans\[3\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13233__CLK clknet_leaf_285_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12914_ _00793_ clknet_leaf_157_clock u2.mem\[49\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06155__A1 u2.mem\[174\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06155__B2 u2.mem\[155\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13383__CLK clknet_leaf_301_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12845_ _00724_ clknet_leaf_205_clock u2.mem\[45\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12776_ _00655_ clknet_leaf_130_clock u2.mem\[40\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07104__B1 _02582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07655__A1 u2.mem\[14\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11727_ _03674_ _05835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07655__B2 u2.mem\[12\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11658_ _05670_ _05792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10609_ _05103_ u2.mem\[58\]\[4\] _05136_ _05137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11589_ _05746_ u2.mem\[174\]\[0\] _05748_ _05749_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13328_ _01207_ clknet_leaf_3_clock u2.mem\[158\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08207__I0 _03554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06091__C2 u2.mem\[161\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13259_ _01138_ clknet_leaf_311_clock u2.mem\[146\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_1546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07820_ u2.mem\[61\]\[12\] _03132_ _03133_ u2.mem\[63\]\[12\] _03287_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07751_ u2.mem\[44\]\[11\] _03120_ _03121_ u2.mem\[42\]\[11\] _03219_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06702_ _02100_ _02186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07682_ _03148_ _03149_ _03150_ _03151_ _03152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06146__A1 _01607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09421_ _04362_ u2.mem\[30\]\[2\] _04396_ _04399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08930__I1 u2.mem\[19\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06633_ u2.mem\[144\]\[0\] _02115_ _02117_ u2.mem\[182\]\[0\] _02118_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07894__A1 u2.mem\[9\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10739__S _05214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12750__CLK clknet_leaf_213_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09352_ _04278_ u2.mem\[28\]\[12\] _04351_ _04352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06564_ _02021_ _02040_ _02048_ _02049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11817__I1 u2.mem\[188\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08209__S _03614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08303_ _03678_ _00086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06449__A2 _01938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08694__I0 _03932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09283_ _04310_ _04311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_166_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06495_ u2.mem\[192\]\[15\] _01981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08234_ _03629_ _03630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_165_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13106__CLK clknet_leaf_241_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08165_ _03589_ _00037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10474__S _05051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07847__I _02602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_241_clock clknet_5_19_0_clock clknet_leaf_241_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_147_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07116_ _02577_ _02578_ _02468_ _02551_ _02595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__07949__A2 _03411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08071__A1 _01958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08096_ _03484_ _03540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12130__CLK clknet_leaf_35_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07047_ _02525_ _02526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06621__A2 _02103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13256__CLK clknet_leaf_311_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_256_clock clknet_5_23_0_clock clknet_leaf_256_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_47_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08998_ _03987_ _04122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12280__CLK clknet_leaf_120_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07949_ _03410_ _03411_ _03412_ _03413_ _03414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_21_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11505__I0 _05677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06198__I _01704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10960_ _03751_ _05354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_95_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09619_ _04498_ u2.mem\[34\]\[15\] _04516_ _04520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10891_ _04072_ _05276_ _05309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_55_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12630_ _00509_ clknet_leaf_96_clock u2.mem\[31\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08119__S _03555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11808__I1 u2.mem\[187\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11998__CLK clknet_leaf_28_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12561_ _00440_ clknet_leaf_170_clock u2.mem\[27\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11512_ _05701_ _01272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10492__I0 _05014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12492_ _00371_ clknet_leaf_190_clock u2.mem\[23\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11443_ _05656_ _01248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_209_clock clknet_5_29_0_clock clknet_leaf_209_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11197__A1 _04179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10244__I0 _04909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06661__I _02145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08062__A1 _03515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11374_ _05613_ _01222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13113_ _00992_ clknet_leaf_327_clock u2.mem\[61\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10325_ _04911_ u2.mem\[51\]\[11\] _04954_ _04958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08789__S _03990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13044_ _00923_ clknet_leaf_26_clock u2.mem\[57\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12623__CLK clknet_leaf_172_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10256_ _04611_ _04918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10187_ _04797_ u2.mem\[48\]\[6\] _04870_ _04873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10172__A2 _04863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12050__D data_in_trans\[0\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06128__A1 _01552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12828_ _00707_ clknet_leaf_208_clock u2.mem\[44\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13129__CLK clknet_leaf_327_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07628__A1 _01954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12759_ _00638_ clknet_leaf_50_clock u2.mem\[39\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10483__I0 _05005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06280_ u2.mem\[187\]\[2\] _01633_ _01636_ u2.mem\[192\]\[2\] _01785_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06300__A1 u2.mem\[147\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06300__B2 u2.mem\[169\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12153__CLK clknet_leaf_56_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13279__CLK clknet_leaf_361_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06851__A2 _02145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08053__A1 _01844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09970_ _04741_ _00690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06603__A2 _02080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08921_ _04017_ u2.mem\[19\]\[1\] _04074_ _04076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09928__I0 _04716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11735__I0 _05825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08852_ _03692_ _04032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_133_clock_I clknet_5_12_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06367__B2 u2.mem\[156\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07803_ u2.mem\[50\]\[12\] _03111_ _03112_ u2.mem\[51\]\[12\] _03270_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08783_ _03984_ _03985_ _03478_ _03986_ _03987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_05995_ _01503_ _01504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07734_ _01962_ _03013_ _03181_ _03202_ _01487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06119__A1 u2.mem\[184\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07867__A1 u2.mem\[32\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07665_ u2.mem\[60\]\[9\] _03055_ _03056_ u2.mem\[62\]\[9\] _03135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11652__I _05787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09404_ _04170_ _04387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06616_ _01992_ _02002_ _02101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07596_ _02569_ _03067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09335_ _04342_ _00454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06547_ _01985_ _02025_ _02032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10474__I0 _04992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09266_ _04301_ _00426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06478_ u2.mem\[193\]\[11\] _01960_ _01948_ u2.mem\[192\]\[11\] _01964_ _01968_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_166_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_180_clock clknet_5_30_0_clock clknet_leaf_180_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08217_ _03620_ _00058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09197_ _04255_ _00403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_58_clock_I clknet_5_12_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09993__S _04750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08148_ _03577_ u2.mem\[1\]\[14\] _03573_ _03578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10932__S _05326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08079_ data_in_trans\[12\].data_sync _03528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_195_clock clknet_5_31_0_clock clknet_leaf_195_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10110_ _04797_ u2.mem\[46\]\[6\] _04825_ _04828_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09919__I0 _04709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11090_ _05420_ u2.mem\[143\]\[0\] _05435_ _05436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09395__I1 u2.mem\[29\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10041_ _04781_ _00721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12796__CLK clknet_leaf_220_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10731__I _03683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06358__B2 u2.mem\[161\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06373__A4 _01875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12026__CLK clknet_leaf_302_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11992_ _00004_ clknet_leaf_329_clock u2.mem\[0\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10943_ _05341_ _01063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_133_clock clknet_5_12_0_clock clknet_leaf_133_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_16_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10874_ _05294_ u2.mem\[130\]\[0\] _05297_ _05298_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_335_clock_I clknet_5_5_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12613_ _00492_ clknet_leaf_94_clock u2.mem\[30\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12176__CLK clknet_leaf_226_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08658__I0 _03908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12544_ _00423_ clknet_leaf_168_clock u2.mem\[26\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_148_clock clknet_5_24_0_clock clknet_leaf_148_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_8_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12475_ _00354_ clknet_leaf_182_clock u2.mem\[22\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06833__A2 _02042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11426_ _04094_ _05645_ _05646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08035__A1 _01545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13571__CLK clknet_leaf_20_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11357_ _05593_ u2.mem\[159\]\[4\] _05597_ _05603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10308_ _04948_ _00821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08312__S _03677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11288_ _05548_ u2.mem\[155\]\[1\] _05559_ _05561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13027_ _00906_ clknet_leaf_42_clock u2.mem\[56\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10239_ _04906_ _00794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06349__A1 u2.mem\[184\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11193__I1 u2.mem\[149\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08111__I _03503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09143__S _04218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11472__I _03506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07450_ u2.mem\[8\]\[5\] _02858_ _02859_ u2.mem\[4\]\[5\] _02924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08982__S _04107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07864__A4 _03330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06401_ u2.mem\[173\]\[5\] _01719_ _01721_ u2.mem\[185\]\[5\] _01903_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07381_ _02618_ _02856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09120_ _04202_ _04208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_52_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06332_ u2.mem\[170\]\[3\] _01687_ _01689_ u2.mem\[156\]\[3\] _01836_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12669__CLK clknet_leaf_193_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09051_ _04163_ _04164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06285__C2 _01645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06263_ u2.mem\[0\]\[2\] _01768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08002_ u2.active_mem\[11\] _03461_ _03462_ u2.active_mem\[10\] _03465_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_102_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06194_ _01700_ _01701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06007__S _01510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11848__S _05905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06588__A1 u2.mem\[184\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09953_ _04731_ _00683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08222__S _03619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08904_ _04039_ u2.mem\[18\]\[11\] _04061_ _04065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12049__CLK clknet_2_3__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09884_ _04686_ _00659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_284_clock_I clknet_5_21_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_11_0_clock clknet_3_5_0_clock clknet_4_11_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_4119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08021__I mem_address_trans\[0\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08835_ _04020_ _00276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08766_ _03928_ u2.mem\[15\]\[10\] _03973_ _03976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07860__I _02621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_50_clock clknet_5_13_0_clock clknet_leaf_50_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_input11_I data_in_a[13] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06760__A1 u2.mem\[188\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07717_ _03182_ _03183_ _03184_ _03185_ _03186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08697_ _03935_ u2.mem\[13\]\[13\] _03933_ _03936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11636__A2 _05769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13444__CLK clknet_leaf_349_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10695__I0 _05115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07648_ u2.mem\[58\]\[9\] _03042_ _03043_ u2.mem\[36\]\[9\] _03118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07579_ _02516_ _03050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_65_clock clknet_5_9_0_clock clknet_leaf_65_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_9_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09318_ _04331_ _00448_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09301__I1 u2.mem\[27\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10590_ _05124_ u2.mem\[57\]\[13\] _05122_ _05125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09249_ _04254_ u2.mem\[26\]\[1\] _04290_ _04292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06276__C2 u2.mem\[176\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12260_ _00139_ clknet_leaf_70_clock u2.mem\[8\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09065__I0 _04174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11211_ _05511_ u2.mem\[150\]\[3\] _05502_ _05512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11758__S _05848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09765__A1 _04180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12191_ _00070_ clknet_leaf_237_clock u2.mem\[4\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11572__A1 _05411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09228__S _04270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput43 net43 driver_io[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_11142_ _05467_ _01136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08132__S _03564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07240__A2 _02546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11557__I _05605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10461__I _05029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11073_ _05339_ _05424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10024_ _04761_ _04772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11875__A2 _05926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08866__I _04014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_18_clock clknet_5_2_0_clock clknet_leaf_18_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06751__A1 u2.mem\[179\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06751__B2 u2.mem\[191\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11975_ _05970_ _05985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_75_1506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10686__I0 _05106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10926_ _05301_ u2.mem\[133\]\[2\] _05327_ _05330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12811__CLK clknet_leaf_221_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10857_ _05286_ _05287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_13_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08307__S _03677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13576_ _01455_ clknet_leaf_32_clock u2.mem\[194\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10788_ _05245_ _01004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12527_ _00406_ clknet_leaf_169_clock u2.mem\[25\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10636__I _05151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12961__CLK clknet_leaf_157_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12458_ _00337_ clknet_leaf_127_clock u2.mem\[20\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07010__I _02488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11668__S _05787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11409_ _05635_ u2.mem\[162\]\[5\] _05624_ _05636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12389_ _00268_ clknet_leaf_78_clock u2.mem\[16\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07767__B1 _03147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07231__A2 _02495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13317__CLK clknet_leaf_301_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06950_ _02362_ _02429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_113_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input3_I col_select_a[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06881_ _02359_ _02360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08620_ _03884_ _00197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13467__CLK clknet_leaf_346_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08551_ _03844_ _00168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07502_ _02970_ _02971_ _02972_ _02973_ _02974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10677__I0 _05097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08482_ _03656_ _03798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07298__A2 _02687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12491__CLK clknet_leaf_182_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09601__S _04506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07433_ _02574_ _02907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07364_ _02584_ _02839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09295__I0 _04260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09103_ _04198_ _00366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09400__I _04166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06315_ _01815_ _01816_ _01817_ _01818_ _01819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_164_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06258__C2 _01653_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07295_ u2.mem\[52\]\[3\] _02601_ _02603_ u2.mem\[21\]\[3\] _02771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09034_ _04150_ _04151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08016__I mem_address_trans\[4\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06246_ u2.mem\[159\]\[1\] _01604_ _01595_ u2.mem\[149\]\[1\] _01752_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07470__A2 _02887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11578__S _05739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06177_ _01683_ _01684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07855__I _02618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07758__B1 _03056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09048__S _04155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10281__I _04922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06430__B1 _01929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09936_ _04687_ u2.mem\[42\]\[2\] _04719_ _04722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09867_ _04675_ _00653_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08686__I _03701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08818_ _03937_ u2.mem\[16\]\[14\] _04005_ _04008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09798_ _04612_ u2.mem\[38\]\[14\] _04633_ _04636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07590__I _02553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06733__A1 u2.mem\[188\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07930__B1 _02561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12834__CLK clknet_leaf_145_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08749_ _03966_ _00244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10668__I0 _05126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11760_ _05837_ u2.mem\[184\]\[5\] _05848_ _05855_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07289__A2 _02565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10711_ _03904_ _05172_ _05195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_1857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10657__S _05162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11691_ _05792_ u2.mem\[180\]\[2\] _05810_ _05813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_1501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12984__CLK clknet_leaf_329_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08238__A1 _03630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13430_ _01309_ clknet_5_4_0_clock u2.mem\[175\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10642_ _05155_ _00948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09286__I0 _04246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06934__I _02412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_23_0_clock_I clknet_4_11_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13361_ _01240_ clknet_leaf_355_clock u2.mem\[163\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10573_ _05094_ _05113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_139_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07997__B1 _03459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12312_ _00191_ clknet_leaf_121_clock u2.mem\[11\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12214__CLK clknet_leaf_68_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13292_ _01171_ clknet_leaf_0_clock u2.mem\[152\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11488__S _05683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12243_ _00122_ clknet_leaf_73_clock u2.mem\[7\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12174_ _00053_ clknet_leaf_210_clock u2.mem\[3\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07213__A2 _02612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12364__CLK clknet_leaf_206_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10191__I _04864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11125_ _05456_ _01130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11056_ _05380_ u2.mem\[141\]\[0\] _05413_ _05414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10007_ _04681_ u2.mem\[44\]\[0\] _04762_ _04763_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06724__A1 u2.mem\[171\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06724__B2 u2.mem\[157\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10659__I0 _05117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11958_ _05909_ u2.mem\[194\]\[2\] _05975_ _05976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09421__S _04396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07819__A4 _03285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10909_ _05320_ _01050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11889_ u2.mem\[192\]\[5\] _03511_ _05932_ _05936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_232_clock_I clknet_5_24_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13559_ _01438_ clknet_leaf_33_clock u2.mem\[193\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07988__B1 _02629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06100_ _01600_ _01607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10831__I0 u2.mem\[63\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07080_ _02558_ _02559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06031_ _01531_ _01534_ _01539_ _01516_ _01540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_160_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12707__CLK clknet_leaf_30_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11387__I1 u2.mem\[161\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07204__A2 _02680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07982_ _03442_ _03443_ _03444_ _03445_ _03446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_86_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06963__A1 _02440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12857__CLK clknet_leaf_133_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06933_ _02346_ _02412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09721_ _04583_ u2.mem\[37\]\[5\] _04580_ _04584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09652_ _04494_ u2.mem\[35\]\[13\] _04537_ _04539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06864_ _01984_ _02008_ _02010_ row_select_trans\[1\].data_sync _02343_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08603_ _03829_ u2.mem\[11\]\[13\] _03872_ _03874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09583_ _04499_ _00545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06795_ u2.mem\[149\]\[4\] _02176_ _02177_ u2.mem\[175\]\[4\] _02276_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06191__A2 _01665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08534_ _03834_ _00161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09331__S _04336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08465_ _03693_ u2.mem\[8\]\[8\] _03788_ _03789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07416_ _02525_ _02890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12237__CLK clknet_leaf_211_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08396_ _03719_ u2.mem\[6\]\[14\] _03743_ _03746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07691__A2 _03013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07347_ _02545_ _02822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07278_ u2.mem\[14\]\[3\] _02657_ _02658_ u2.mem\[12\]\[3\] _02754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_128_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09017_ _04137_ _00341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12387__CLK clknet_leaf_77_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06229_ u2.mem\[145\]\[1\] _01640_ _01734_ u2.mem\[177\]\[1\] _01735_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07585__I _02548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06403__B1 _01683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09919_ _04709_ u2.mem\[41\]\[12\] _04710_ _04711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_181_clock_I clknet_5_30_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12930_ _00809_ clknet_leaf_234_clock u2.mem\[50\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10889__I0 _05307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06929__I _02389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06706__A1 _02184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12861_ _00740_ clknet_leaf_200_clock u2.mem\[46\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13012__CLK clknet_leaf_31_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11812_ _05887_ _05888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12792_ _00671_ clknet_leaf_44_clock u2.mem\[41\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11743_ _05835_ u2.mem\[183\]\[4\] _05839_ _05845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11674_ _05790_ u2.mem\[179\]\[1\] _05801_ _05803_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13162__CLK clknet_leaf_275_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11066__I0 _05392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13413_ _01292_ clknet_leaf_344_clock u2.mem\[172\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10625_ _05145_ _00941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07434__A2 _02906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13344_ _01223_ clknet_leaf_8_clock u2.mem\[160\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10556_ _04997_ _05101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13275_ _01154_ clknet_leaf_12_clock u2.mem\[149\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10487_ _05009_ u2.mem\[55\]\[7\] _05056_ _05060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11369__I1 u2.mem\[160\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12226_ _00105_ clknet_leaf_143_clock u2.mem\[6\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07198__A1 u2.mem\[29\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11946__S _05965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12157_ _00036_ clknet_leaf_205_clock u2.mem\[2\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12053__D net15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11108_ _05424_ u2.mem\[144\]\[1\] _05445_ _05447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12088_ row_col_select_trans.A clknet_leaf_298_clock row_col_select_trans.data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09734__I1 u2.mem\[37\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11039_ _04334_ _05402_ _05403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_37_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06580_ _02064_ _02028_ _02065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09498__I0 _04360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09151__S _04226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13505__CLK clknet_leaf_318_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10297__S _04938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08250_ _03641_ _00070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07673__A2 _03069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07201_ _02675_ _02676_ _02677_ _02678_ _02679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_105_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08181_ _03598_ _00044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10096__I _04819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07132_ _02566_ _02567_ _02404_ _02568_ _02611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__09670__I0 _04473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07063_ _02541_ _02542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11509__A1 _04248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06014_ u2.driver_mem\[7\] _01508_ _01523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_138_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08225__I1 u2.mem\[3\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07965_ u2.mem\[58\]\[15\] _03275_ _03276_ u2.mem\[36\]\[15\] _03429_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11655__I _05667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13035__CLK clknet_leaf_248_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09704_ _04570_ u2.mem\[37\]\[1\] _04567_ _04571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06916_ _02388_ _02390_ _02393_ _02394_ _02395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_60_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07896_ _03358_ _03359_ _03360_ _03361_ _03362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_112_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11532__I1 u2.mem\[170\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09635_ _04529_ _00567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06847_ u2.mem\[148\]\[5\] _02128_ _02130_ u2.mem\[152\]\[5\] _02327_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09489__I0 _04391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09566_ _04487_ u2.mem\[33\]\[10\] _04483_ _04488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06778_ _02256_ _02257_ _02258_ _02259_ _02260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_55_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08517_ _03822_ u2.mem\[9\]\[10\] _03818_ _03823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11296__I0 _05556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09497_ _04444_ _00514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09996__S _04755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10000__S _04755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08448_ _03779_ _00130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07664__A2 _03132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_128_clock_I clknet_5_14_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08379_ _03736_ _00104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11748__A1 _04223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10410_ _05013_ _00858_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11390_ _05622_ _01229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09661__I0 _04463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10341_ _04889_ u2.mem\[52\]\[1\] _04966_ _04968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10734__I _03687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13060_ _00939_ clknet_leaf_27_clock u2.mem\[58\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10272_ _04922_ _04928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_65_1313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12011_ net27 clknet_2_1__leaf_clock_a mem_address_trans\[3\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11766__S _05857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06659__I _02143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12402__CLK clknet_leaf_155_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13528__CLK clknet_leaf_317_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12913_ _00792_ clknet_leaf_158_clock u2.mem\[49\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12844_ _00723_ clknet_leaf_204_clock u2.mem\[45\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12775_ _00654_ clknet_leaf_131_clock u2.mem\[40\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12552__CLK clknet_leaf_119_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11726_ _05834_ _01353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07655__A2 _03123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06312__C1 _01660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11657_ _05791_ _01327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10845__S _05278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10608_ _05130_ _05136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_167_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09652__I0 _04494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11588_ _05747_ _05748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_143_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13327_ _01206_ clknet_leaf_3_clock u2.mem\[158\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10539_ _05023_ u2.mem\[56\]\[13\] _05088_ _05090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06091__B2 u2.mem\[149\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08114__I _03507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13258_ _01137_ clknet_leaf_312_clock u2.mem\[146\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11676__S _05801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13058__CLK clknet_leaf_242_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12209_ _00088_ clknet_leaf_232_clock u2.mem\[5\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10580__S _05113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_1574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13189_ _01068_ clknet_leaf_277_clock u2.mem\[135\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06918__B2 u2.mem\[2\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11911__A1 _03535_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06394__A2 _01889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07750_ _03214_ _03215_ _03216_ _03217_ _03218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_133_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12082__CLK clknet_leaf_363_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06701_ _02103_ _02185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07681_ u2.mem\[18\]\[9\] _03083_ _03084_ u2.mem\[19\]\[9\] _03151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06146__A2 _01629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07343__B2 u2.mem\[20\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09420_ _04398_ _00483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06632_ _02116_ _02117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08784__I _03987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09351_ _04335_ _04351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06563_ u2.mem\[180\]\[0\] _02043_ _02047_ u2.mem\[150\]\[0\] _02048_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10819__I _05252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08302_ _03676_ u2.mem\[5\]\[4\] _03677_ _03678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09282_ _03748_ _04247_ _04310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06494_ u2.mem\[0\]\[15\] _01980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07646__A2 _03114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08233_ mem_address_trans\[1\].data_sync mem_address_trans\[0\].data_sync _03629_
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_165_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08164_ _03552_ u2.mem\[2\]\[3\] _03585_ _03589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09643__I0 _04485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07115_ u2.mem\[17\]\[0\] _02591_ _02593_ u2.mem\[24\]\[0\] _02594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_174_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07949__A3 _03412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11450__I0 _05633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08095_ _03492_ _03539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08071__A2 _03517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06082__A1 _01586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07046_ _02466_ _02467_ _02411_ _02394_ _02525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_162_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10490__S _05061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input41_I row_select_a[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12425__CLK clknet_leaf_128_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06385__A2 _01884_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08997_ _04120_ _04121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07582__A1 _03024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07948_ u2.mem\[6\]\[14\] _03327_ _03328_ u2.mem\[47\]\[14\] _03413_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_5_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_54_clock_I clknet_5_12_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11505__I1 u2.mem\[168\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09323__A2 _04334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07879_ u2.mem\[58\]\[13\] _03275_ _03276_ u2.mem\[36\]\[13\] _03345_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12575__CLK clknet_leaf_183_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09618_ _04519_ _00560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10890_ _05308_ _01043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09549_ _04144_ _04476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12560_ _00439_ clknet_leaf_171_clock u2.mem\[27\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07637__A2 _03028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07103__I _02581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06845__B1 _02134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11511_ _05663_ u2.mem\[169\]\[0\] _05700_ _05701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_279_clock_I clknet_5_21_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12491_ _00370_ clknet_leaf_182_clock u2.mem\[23\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06942__I _02402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11442_ _05623_ u2.mem\[165\]\[0\] _05655_ _05656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09634__I0 _04476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08135__S _03564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11197__A2 _05482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11373_ _05593_ u2.mem\[160\]\[4\] _05607_ _05613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13200__CLK clknet_leaf_271_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10324_ _04957_ _00828_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13112_ _00991_ clknet_leaf_39_clock u2.mem\[61\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_331_clock_I clknet_5_7_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10255_ _04917_ _00799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13043_ _00922_ clknet_leaf_26_clock u2.mem\[57\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_363_clock clknet_5_0_0_clock clknet_leaf_363_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08869__I _03714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10186_ _04872_ _00775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12918__CLK clknet_leaf_84_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06781__C1 u2.mem\[181\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06128__A2 _01634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10180__I0 _04790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07876__A2 _02503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12827_ _00706_ clknet_leaf_221_clock u2.mem\[44\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_301_clock clknet_5_16_0_clock clknet_leaf_301_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_61_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08125__I0 _03561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07628__A2 _03013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12758_ _00637_ clknet_leaf_74_clock u2.mem\[39\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09873__I0 _04612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07013__I _02432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11680__I0 _05796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11709_ _05796_ u2.mem\[181\]\[4\] _05817_ _05823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06836__B1 _02105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12689_ _00568_ clknet_leaf_174_clock u2.mem\[35\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06300__A2 _01676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_316_clock clknet_5_18_0_clock clknet_leaf_316_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_163_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09625__I0 _04467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11432__I0 _05629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10374__I _04117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06064__A1 _01547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12448__CLK clknet_leaf_159_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07261__B1 _02634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08920_ _04075_ _00306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07683__I _02626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11735__I1 u2.mem\[183\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08851_ _04031_ _00281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06367__A2 _01686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12598__CLK clknet_leaf_96_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07802_ _03260_ _03263_ _03266_ _03268_ _03269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06906__A4 _02384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08782_ mem_address_trans\[7\].data_sync _03986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05994_ u2.select_mem_row\[1\] u2.select_mem_col\[1\] _01502_ _01503_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09604__S _04511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07733_ _03186_ _03191_ _03196_ _03201_ _03202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__11499__I0 _05668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07664_ u2.mem\[61\]\[9\] _03132_ _03133_ u2.mem\[63\]\[9\] _03134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09403_ _04386_ _00478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06615_ _02028_ _02053_ _02100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_164_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07595_ _02564_ _03066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08116__I0 _03554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09334_ _04260_ u2.mem\[28\]\[4\] _04341_ _04342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06546_ _02006_ _02031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07619__A2 _03088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08019__I _03479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09864__I0 _04599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_280_clock_I clknet_5_21_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09265_ _04269_ u2.mem\[26\]\[8\] _04300_ _04301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06477_ u2.mem\[194\]\[11\] _01946_ _01967_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10485__S _05056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13223__CLK clknet_leaf_286_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07858__I _02613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08216_ _03563_ u2.mem\[3\]\[8\] _03619_ _03620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09196_ _04254_ u2.mem\[25\]\[1\] _04252_ _04255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11423__I0 _05635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08147_ _03533_ _03577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07252__B1 _02608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08078_ _03489_ _03527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13373__CLK clknet_leaf_354_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07029_ _02413_ _02491_ _02492_ _02507_ _02508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_136_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08689__I _03705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10040_ _04716_ u2.mem\[44\]\[15\] _04777_ _04781_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06430__C _01914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09514__S _04453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11991_ _00003_ clknet_leaf_318_clock u2.mem\[0\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10942_ _05340_ u2.mem\[134\]\[1\] _05337_ _05341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10873_ _05296_ _05297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_12612_ _00491_ clknet_leaf_93_clock u2.mem\[30\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09855__I0 _04586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12543_ _00422_ clknet_leaf_168_clock u2.mem\[26\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11662__I0 _05794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10395__S _05002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06294__A1 u2.mem\[144\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07491__B1 _02921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06294__B2 u2.mem\[182\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12474_ _00353_ clknet_leaf_123_clock u2.mem\[21\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11425_ _05605_ _05645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_158_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06046__A1 _01547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11356_ _05602_ _01215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10307_ _04893_ u2.mem\[51\]\[3\] _04944_ _04948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12740__CLK clknet_leaf_67_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11287_ _05560_ _01188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13026_ _00905_ clknet_leaf_251_clock u2.mem\[56\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10238_ _04904_ u2.mem\[49\]\[8\] _04905_ _04906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07546__A1 u2.mem\[32\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08594__I0 _03820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07546__B2 u2.mem\[2\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12061__D net19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10169_ _03477_ mem_address_trans\[5\].data_sync _04861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07008__I _02346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12890__CLK clknet_leaf_140_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_240_clock clknet_5_19_0_clock clknet_leaf_240_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_130_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13246__CLK clknet_leaf_272_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06400_ u2.mem\[144\]\[5\] _01670_ _01672_ u2.mem\[182\]\[5\] _01902_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06521__A2 row_select_trans\[4\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07380_ _02616_ _02855_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09846__I0 _04573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06331_ u2.mem\[173\]\[3\] _01720_ _01722_ u2.mem\[185\]\[3\] _01835_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_255_clock clknet_5_23_0_clock clknet_leaf_255_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11653__I0 _05786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09050_ data_in_trans\[11\].data_sync _04163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06285__A1 u2.mem\[145\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06285__B2 u2.mem\[163\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06262_ _01727_ _01554_ _01737_ _01767_ _01481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12270__CLK clknet_leaf_185_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08001_ _03460_ _03463_ _03464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06193_ _01615_ _01596_ _01700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07234__B1 _02658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09952_ _04703_ u2.mem\[42\]\[9\] _04729_ _04731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08903_ _04064_ _00300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09883_ _04685_ u2.mem\[41\]\[1\] _04683_ _04686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_227_clock_I clknet_5_25_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08585__I0 _03811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08834_ _04019_ u2.mem\[17\]\[2\] _04015_ _04020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08765_ _03975_ _00251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_208_clock clknet_5_29_0_clock clknet_leaf_208_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_96_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07716_ u2.mem\[57\]\[10\] _03061_ _03062_ u2.mem\[41\]\[10\] _03185_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08696_ _03714_ _03935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07647_ u2.mem\[53\]\[9\] _03039_ _03040_ u2.mem\[56\]\[9\] _03117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_14_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07578_ _02514_ _03049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09837__I0 _04615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12613__CLK clknet_leaf_94_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09317_ _04283_ u2.mem\[27\]\[14\] _04328_ _04331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06529_ _02013_ _02014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11644__I0 _05754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07588__I _02541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06276__A1 u2.mem\[189\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09248_ _04291_ _00418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06276__B2 u2.mem\[180\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09179_ _04242_ _00398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12763__CLK clknet_leaf_203_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07225__B1 _02477_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11210_ _05510_ _05511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12190_ _00069_ clknet_leaf_252_clock u2.mem\[4\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11572__A2 _05729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11141_ _05466_ u2.mem\[146\]\[2\] _05462_ _05467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput44 net44 driver_io[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_1_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13119__CLK clknet_leaf_243_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11072_ _05423_ _01110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08576__I0 _03802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10023_ _04771_ _00713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06200__A1 _01556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12143__CLK clknet_leaf_218_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08328__I0 _03698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11573__I _05738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13269__CLK clknet_leaf_5_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06751__A2 _02150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11088__A1 _04417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11974_ _05984_ _01451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09043__I _04157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10925_ _05329_ _01057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11883__I0 u2.mem\[192\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12293__CLK clknet_leaf_101_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09828__I0 _04602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10856_ _05285_ _05276_ _05286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_60_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_13575_ _01454_ clknet_leaf_34_clock u2.mem\[194\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10787_ _05218_ u2.mem\[62\]\[10\] _05242_ _05245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12526_ _00405_ clknet_leaf_187_clock u2.mem\[25\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12056__D data_in_trans\[3\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12457_ _00336_ clknet_leaf_126_clock u2.mem\[20\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10853__S _05277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09419__S _04396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11408_ _05516_ _05635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06019__B2 _01516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08323__S _03694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12388_ _00267_ clknet_leaf_81_clock u2.mem\[16\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11339_ _05591_ u2.mem\[158\]\[3\] _05585_ _05592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09218__I _04251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07519__A1 _02974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13009_ _00888_ clknet_leaf_239_clock u2.mem\[55\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06880_ _02358_ _02359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07534__A4 _03005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08550_ _03813_ u2.mem\[10\]\[6\] _03841_ _03844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10126__I0 _04813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12636__CLK clknet_leaf_192_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07501_ u2.mem\[27\]\[7\] _02788_ _02789_ u2.mem\[35\]\[7\] _02973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08481_ _03797_ _00145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07432_ _02572_ _02906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_194_clock clknet_5_31_0_clock clknet_leaf_194_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09819__I0 _04589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11626__I0 _05750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07363_ u2.mem\[9\]\[4\] _02836_ _02837_ u2.mem\[25\]\[4\] _02838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09295__I1 u2.mem\[27\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12786__CLK clknet_leaf_321_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09102_ _04167_ u2.mem\[22\]\[12\] _04197_ _04198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06258__A1 u2.mem\[189\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07455__B1 _02867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06314_ u2.mem\[172\]\[3\] _01654_ _01664_ u2.mem\[180\]\[3\] _01818_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06258__B2 u2.mem\[176\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07294_ u2.mem\[17\]\[3\] _02591_ _02593_ u2.mem\[24\]\[3\] _02770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09033_ data_in_trans\[7\].data_sync _04150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06245_ _01746_ _01747_ _01748_ _01750_ _01751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_164_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09329__S _04336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07207__B1 _02608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06176_ _01581_ _01641_ _01683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_132_clock clknet_5_12_0_clock clknet_leaf_132_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_131_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06430__A1 u2.mem\[193\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09935_ _04721_ _00675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06430__B2 u2.mem\[192\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08032__I _03488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12166__CLK clknet_leaf_91_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09866_ _04602_ u2.mem\[40\]\[11\] _04671_ _04675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13411__CLK clknet_leaf_341_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06718__C1 _02019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_147_clock clknet_5_24_0_clock clknet_leaf_147_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08817_ _04007_ _00271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09797_ _04635_ _00623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11393__I _05624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10117__I0 _04804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08748_ _03910_ u2.mem\[15\]\[2\] _03963_ _03966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13561__CLK clknet_leaf_32_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11865__I0 _05909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08679_ _03692_ _03923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10938__S _05337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_9_0_clock clknet_3_4_0_clock clknet_4_9_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_41_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10710_ _04986_ _05194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11690_ _05812_ _01339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10641_ _05099_ u2.mem\[59\]\[2\] _05152_ _05155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10737__I _03691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09286__I1 u2.mem\[27\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13360_ _01239_ clknet_leaf_356_clock u2.mem\[163\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06249__B2 u2.mem\[161\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10572_ _03691_ _05112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12311_ _00190_ clknet_leaf_118_clock u2.mem\[11\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13291_ _01170_ clknet_leaf_361_clock u2.mem\[152\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_5_27_0_clock_I clknet_4_13_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06950__I _02362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12242_ _00121_ clknet_leaf_226_clock u2.mem\[7\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07749__B2 u2.mem\[36\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12509__CLK clknet_leaf_180_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12173_ _00052_ clknet_leaf_210_clock u2.mem\[3\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09038__I _04153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11124_ _05426_ u2.mem\[145\]\[2\] _05453_ _05456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13091__CLK clknet_leaf_22_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11055_ _05412_ _05413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07781__I _02385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10006_ _04761_ _04762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_77_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07921__A1 u2.mem\[53\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07921__B2 u2.mem\[56\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10108__I0 _04795_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11957_ _05971_ _05975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_79_1495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06488__A1 _01973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07685__B1 _03154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10908_ _05294_ u2.mem\[132\]\[0\] _05319_ _05320_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11888_ _05935_ _01414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11608__I0 _05746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10839_ _03477_ _03985_ _05274_ _05275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_38_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12039__CLK clknet_2_2__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13558_ _01437_ clknet_leaf_19_clock u2.mem\[193\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07021__I _02499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12509_ _00388_ clknet_leaf_180_clock u2.mem\[24\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10583__S _05113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10831__I1 _03531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07452__A3 _02924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13489_ _01368_ clknet_leaf_293_clock u2.mem\[185\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06030_ _01504_ _01536_ _01538_ _01539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12189__CLK clknet_leaf_252_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06412__A1 _01911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07981_ u2.mem\[28\]\[15\] _03305_ _03306_ u2.mem\[31\]\[15\] _03445_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_45_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_64_clock clknet_5_9_0_clock clknet_leaf_64_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06963__A2 _02441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09720_ _04582_ _04583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06932_ _02410_ _02403_ _02392_ _02411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_67_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09651_ _04538_ _00574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06863_ col_select_trans\[5\].data_sync _02024_ _02016_ col_select_trans\[4\].data_sync
+ _02342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_82_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07912__A1 u2.mem\[27\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08602_ _03873_ _00190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08960__I0 _04017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09582_ _04498_ u2.mem\[33\]\[15\] _04492_ _04499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06794_ u2.mem\[166\]\[4\] _02096_ _02098_ u2.mem\[161\]\[4\] u2.mem\[159\]\[4\]
+ _02174_ _02275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_55_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_79_clock clknet_5_8_0_clock clknet_leaf_79_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_36_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06191__A3 _01678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08533_ _03833_ u2.mem\[9\]\[15\] _03827_ _03834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06100__I _01600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11941__I _05949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06479__A1 _01966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08464_ _03777_ _03788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_24_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07415_ u2.mem\[44\]\[5\] _02887_ _02888_ u2.mem\[42\]\[5\] _02889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08395_ _03745_ _00111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07346_ u2.mem\[61\]\[4\] _02666_ _02667_ u2.mem\[63\]\[4\] _02821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07979__A1 u2.mem\[29\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11589__S _05748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07979__B2 u2.mem\[11\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10822__I1 _03521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07277_ u2.mem\[44\]\[3\] _02654_ _02655_ u2.mem\[42\]\[3\] _02753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_17_clock clknet_5_2_0_clock clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_163_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09016_ _04136_ u2.mem\[21\]\[3\] _04124_ _04137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06228_ _01583_ _01734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06159_ _01638_ _01665_ _01591_ _01666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_144_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08898__S _04061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06403__A1 u2.mem\[191\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07600__B1 _03070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09918_ _04682_ _04710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_63_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08156__A1 _03480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_124_clock_I clknet_5_15_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09849_ _04665_ _00645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06706__A2 _02188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12860_ _00739_ clknet_leaf_203_clock u2.mem\[46\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12951__CLK clknet_leaf_49_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07106__I _02584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11811_ _04333_ _05886_ _05887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_61_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12791_ _00670_ clknet_leaf_44_clock u2.mem\[41\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08703__I0 _03939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11742_ _05844_ _01359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08138__S _03564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10510__I0 _04987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13307__CLK clknet_leaf_359_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11673_ _05802_ _01332_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13412_ _01291_ clknet_leaf_344_clock u2.mem\[172\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10624_ _05119_ u2.mem\[58\]\[11\] _05141_ _05145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11499__S _05692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13343_ _01222_ clknet_leaf_3_clock u2.mem\[160\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12331__CLK clknet_leaf_207_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10813__I1 _03511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10555_ _05100_ _00916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_49_clock_I clknet_5_7_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13457__CLK clknet_leaf_304_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06642__A1 _02007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13274_ _01153_ clknet_leaf_13_clock u2.mem\[149\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10486_ _05059_ _00888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11298__I _05442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12225_ _00104_ clknet_leaf_232_clock u2.mem\[6\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10577__I0 _05115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07198__A2 _02565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12481__CLK clknet_leaf_164_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12156_ _00035_ clknet_leaf_205_clock u2.mem\[2\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08601__S _03872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06945__A2 _02423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11107_ _05446_ _01122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12087_ net36 clknet_2_1__leaf_clock_a row_col_select_trans.A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11038_ _05275_ _05402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_42_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11962__S _05975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07016__I _02494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11829__I0 _05868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09498__I1 u2.mem\[32\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12989_ _00868_ clknet_leaf_258_clock u2.mem\[54\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07658__B1 _03127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10501__I0 _05023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09231__I _04251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_326_clock_I clknet_5_7_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10377__I _04988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06330__B1 _01700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07200_ u2.mem\[28\]\[1\] _02585_ _02587_ u2.mem\[31\]\[1\] _02678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08180_ _03568_ u2.mem\[2\]\[10\] _03595_ _03598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07131_ _02594_ _02599_ _02604_ _02609_ _02610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_146_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10804__I1 _03497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07062_ _02426_ _02399_ _02400_ _02425_ _02541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__06633__A1 u2.mem\[144\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06633__B2 u2.mem\[182\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11509__A2 _05690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06013_ _01516_ _01521_ _01522_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_161_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08511__S _03818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06397__B1 _01714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10840__I _05275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12974__CLK clknet_leaf_261_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07964_ u2.mem\[53\]\[15\] _03272_ _03273_ u2.mem\[56\]\[15\] _03428_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09703_ _04569_ _04570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06915_ _02363_ _02394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08310__I _03683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07895_ u2.mem\[28\]\[13\] _03305_ _03306_ u2.mem\[31\]\[13\] _03361_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09634_ _04476_ u2.mem\[35\]\[5\] _04527_ _04529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07897__B1 _02598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06846_ u2.mem\[153\]\[5\] _02136_ _02137_ u2.mem\[160\]\[5\] _02326_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12204__CLK clknet_leaf_211_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09565_ _04160_ _04487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06777_ u2.mem\[145\]\[3\] _02081_ _02091_ u2.mem\[177\]\[3\] _02259_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_70_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11671__I _05800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08516_ _03701_ _03822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11296__I1 u2.mem\[155\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09496_ _04356_ u2.mem\[32\]\[0\] _04443_ _04444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08447_ _03657_ u2.mem\[8\]\[0\] _03778_ _03779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12354__CLK clknet_leaf_150_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08378_ _03685_ u2.mem\[6\]\[6\] _03733_ _03736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11748__A2 _05847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07329_ u2.mem\[50\]\[4\] _02645_ _02646_ u2.mem\[51\]\[4\] _02804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_50_clock_I clknet_5_13_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07596__I _02569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09661__I1 u2.mem\[36\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11112__S _05445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06624__A1 _02108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10340_ _04967_ _00834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10271_ _04927_ _00805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12010_ mem_address_trans\[2\].A clknet_leaf_312_clock mem_address_trans\[2\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06388__B1 _01732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10750__I _03708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_275_clock_I clknet_5_21_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11782__S _05866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12912_ _00791_ clknet_leaf_147_clock u2.mem\[49\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12843_ _00722_ clknet_leaf_198_clock u2.mem\[45\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12774_ _00653_ clknet_leaf_79_clock u2.mem\[40\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09051__I _04163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07104__A2 _02580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_6_0_clock clknet_0_clock clknet_3_6_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_1463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11987__A2 _05972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11725_ _05833_ u2.mem\[182\]\[3\] _05827_ _05834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06312__B1 _01666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06312__C2 u2.mem\[181\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09986__I _04739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06863__A1 col_select_trans\[5\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11656_ _05790_ u2.mem\[178\]\[1\] _05788_ _05791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12847__CLK clknet_leaf_151_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10607_ _05135_ _00933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11587_ _04393_ _05729_ _05747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_155_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11022__S _05381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10798__I0 _05229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13326_ _01205_ clknet_leaf_304_clock u2.mem\[157\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06615__A1 _02028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07812__B1 _03121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10538_ _05089_ _00910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06091__A2 _01592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13257_ _01136_ clknet_leaf_312_clock u2.mem\[146\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10469_ _05049_ _00881_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12208_ _00087_ clknet_leaf_231_clock u2.mem\[5\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11211__I1 u2.mem\[150\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13188_ _01067_ clknet_leaf_270_clock u2.mem\[134\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07040__A1 _02410_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12139_ _00018_ clknet_leaf_212_clock u2.mem\[1\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12227__CLK clknet_leaf_64_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06700_ u2.mem\[171\]\[1\] _02065_ _02067_ u2.mem\[157\]\[1\] _02183_ _02184_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_07680_ u2.mem\[52\]\[9\] _03080_ _03081_ u2.mem\[21\]\[9\] _03150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10722__I0 _05202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06631_ _02000_ _02046_ _02116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_93_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12377__CLK clknet_leaf_60_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09350_ _04350_ _00461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10101__S _04820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06562_ _02045_ _02046_ _02047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09340__I0 _04267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08301_ _03659_ _03677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_33_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09281_ _04309_ _00433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06493_ u2.mem\[194\]\[15\] _01979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08232_ _03628_ _00065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08163_ _03588_ _00036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10789__I0 _05220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07114_ _02592_ _02593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06606__A1 _02080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07803__B1 _03112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08305__I _03679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08094_ _03537_ _03538_ _00017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11450__I1 u2.mem\[165\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_8_0_clock clknet_4_4_0_clock clknet_5_8_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_88_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07045_ u2.mem\[44\]\[0\] _02521_ _02523_ u2.mem\[42\]\[0\] _02524_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06082__A2 _01588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10771__S _05232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13002__CLK clknet_leaf_322_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07031__A1 _02487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08996_ _03901_ _03750_ _04120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_9_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07582__A2 _03036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input34_I mem_write_n_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13152__CLK clknet_leaf_245_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08040__I data_in_trans\[2\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07947_ u2.mem\[8\]\[14\] _03324_ _03325_ u2.mem\[4\]\[14\] _03412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08975__I _04096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10713__I0 _05194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07878_ u2.mem\[53\]\[13\] _03272_ _03273_ u2.mem\[56\]\[13\] _03344_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09617_ _04496_ u2.mem\[34\]\[14\] _04516_ _04519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06829_ _02305_ _02306_ _02307_ _02308_ _02309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_28_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10011__S _04762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09548_ _04475_ _00534_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09331__I0 _04258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09800__S _04633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09479_ _04432_ _00508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10946__S _05337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11510_ _05699_ _05700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_12_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06845__A1 u2.mem\[194\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12490_ _00369_ clknet_leaf_121_clock u2.mem\[22\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06845__B2 u2.mem\[190\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11441_ _05654_ _05655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08215__I _03608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11372_ _05612_ _01221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13111_ _00990_ clknet_leaf_38_clock u2.mem\[61\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10323_ _04909_ u2.mem\[51\]\[10\] _04954_ _04957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10681__S _05174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09247__S _04290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09398__I0 _04382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13042_ _00921_ clknet_leaf_321_clock u2.mem\[57\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10254_ _04916_ u2.mem\[49\]\[13\] _04914_ _04917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10480__I _05050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07022__B2 u2.mem\[36\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10185_ _04795_ u2.mem\[48\]\[5\] _04870_ _04872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09046__I data_in_trans\[10\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06781__B1 _02034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06781__C2 _02038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10704__I0 _05124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12826_ _00705_ clknet_leaf_136_clock u2.mem\[43\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12059__D net18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12757_ _00636_ clknet_leaf_70_clock u2.mem\[39\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11708_ _05822_ _01347_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06836__A1 u2.mem\[188\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12688_ _00567_ clknet_leaf_177_clock u2.mem\[35\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11680__I1 u2.mem\[179\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13025__CLK clknet_leaf_251_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11639_ _05780_ _01320_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11432__I1 u2.mem\[164\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13309_ _01188_ clknet_leaf_348_clock u2.mem\[155\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06064__A2 _01570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09389__I0 _04375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09157__S _04226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08850_ _04030_ u2.mem\[17\]\[7\] _04024_ _04031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07801_ u2.mem\[3\]\[12\] _03267_ _03211_ _03268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07564__A2 _03034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08781_ mem_address_trans\[5\].data_sync _03985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_22_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05993_ row_col_select_trans.data_sync _01502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07732_ _03197_ _03198_ _03199_ _03200_ _03201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08795__I _03989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07663_ _02560_ _03133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09402_ _04384_ u2.mem\[29\]\[12\] _04385_ _04386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06614_ _02098_ _02099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07594_ u2.mem\[26\]\[8\] _02906_ _02907_ u2.mem\[10\]\[8\] _03065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09313__I0 _04278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09333_ _04335_ _04341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_55_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06545_ _02029_ _02030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11120__I0 _05420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_223_clock_I clknet_5_25_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09264_ _04289_ _04300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06827__B2 u2.mem\[183\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06476_ u2.mem\[0\]\[11\] _01966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08215_ _03608_ _03619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_21_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09195_ _04127_ _04254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08146_ _03576_ _00031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11423__I1 u2.mem\[163\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13518__CLK clknet_leaf_330_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08077_ _01966_ _03517_ _03526_ _00012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07028_ _02441_ _02382_ _02392_ _02507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_162_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11187__I0 _05466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11396__I _05504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12542__CLK clknet_leaf_188_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07095__B _02493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08979_ _04109_ _00331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11990_ _00002_ clknet_leaf_329_clock u2.mem\[0\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10941_ _05339_ _05340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10872_ _05295_ _05276_ _05296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_44_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09304__I0 _04269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07114__I _02592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_12611_ _00490_ clknet_leaf_94_clock u2.mem\[30\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13048__CLK clknet_leaf_44_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09855__I1 u2.mem\[40\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12542_ _00421_ clknet_leaf_188_clock u2.mem\[26\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06953__I _02373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11811__A1 _04333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11662__I1 u2.mem\[178\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12473_ _00352_ clknet_leaf_122_clock u2.mem\[21\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11424_ _05644_ _01241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13198__CLK clknet_leaf_276_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12072__CLK clknet_leaf_28_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06046__A2 _01549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07243__A1 _02716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08291__I0 _03668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11355_ _05591_ u2.mem\[159\]\[3\] _05598_ _05602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07784__I _02405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10306_ _04947_ _00820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11286_ _05544_ u2.mem\[155\]\[0\] _05559_ _05560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13025_ _00904_ clknet_leaf_251_clock u2.mem\[56\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10237_ _04886_ _04905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_105_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09791__I0 _04602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10168_ _04860_ _00769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06754__B1 _02143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_172_clock_I clknet_5_27_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10099_ _04786_ u2.mem\[46\]\[1\] _04820_ _04822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09504__I _04442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09543__I0 _04471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07024__I _02502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12809_ _00688_ clknet_leaf_139_clock u2.mem\[42\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06330_ u2.mem\[154\]\[3\] _01698_ _01700_ u2.mem\[162\]\[3\] _01833_ _01834_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_52_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11653__I1 u2.mem\[178\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06285__A2 _01639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06261_ _01745_ _01751_ _01758_ _01766_ _01767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_31_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10385__I _04994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07482__B2 u2.mem\[11\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08000_ u2.active_mem\[7\] _03461_ _03462_ u2.active_mem\[6\] _03463_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_128_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06192_ _01698_ _01699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_50_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_97_clock_I clknet_5_10_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12565__CLK clknet_leaf_96_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07234__B2 u2.mem\[12\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09951_ _04730_ _00682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11169__I0 _05460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06993__B1 _02471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08902_ _04037_ u2.mem\[18\]\[10\] _04061_ _04064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09882_ _04569_ _04685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10916__I0 _05305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08585__I1 u2.mem\[11\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08833_ _03667_ _04019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09782__I0 _04589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08764_ _03926_ u2.mem\[15\]\[9\] _03973_ _03975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09534__I0 _04463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09414__I _04393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07715_ u2.mem\[37\]\[10\] _03058_ _03059_ u2.mem\[59\]\[10\] _03184_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08695_ _03934_ _00222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_2_3__f_clock_a clknet_0_clock_a clknet_2_3__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_22_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07646_ u2.mem\[54\]\[9\] _03114_ _03115_ u2.mem\[55\]\[9\] _03116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11892__I1 _03513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07577_ u2.mem\[49\]\[8\] _02893_ _02894_ u2.mem\[46\]\[8\] _03048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10496__S _05061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_362_clock clknet_5_0_0_clock clknet_leaf_362_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_41_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09316_ _04330_ _00447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12095__CLK clknet_leaf_214_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06528_ _02007_ _02012_ _02013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13340__CLK clknet_leaf_4_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09247_ _04246_ u2.mem\[26\]\[0\] _04290_ _04291_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07473__B2 u2.mem\[20\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06459_ u2.mem\[193\]\[7\] _01942_ _01948_ u2.mem\[192\]\[7\] _01949_ _01953_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_107_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12908__CLK clknet_leaf_202_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09178_ _04167_ u2.mem\[24\]\[12\] _04241_ _04242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08129_ _03563_ u2.mem\[1\]\[8\] _03564_ _03565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08273__I0 _03579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13490__CLK clknet_leaf_292_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11120__S _05453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10080__I0 _04808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07776__A2 _03241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11140_ _05342_ _05466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_4_5_0_clock clknet_3_2_0_clock clknet_4_5_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_107_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_300_clock clknet_5_17_0_clock clknet_leaf_300_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_1_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11071_ _05420_ u2.mem\[142\]\[0\] _05422_ _05423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09525__S _04458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10022_ _04698_ u2.mem\[44\]\[7\] _04767_ _04771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09773__I0 _04576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11580__I0 _05715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06200__A2 _01677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_315_clock clknet_5_18_0_clock clknet_leaf_315_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09324__I _04335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09525__I0 _04387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11973_ _05216_ u2.mem\[194\]\[9\] _05980_ _05984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10924_ _05299_ u2.mem\[133\]\[1\] _05327_ _05329_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11883__I1 _03500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09260__S _04295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07700__A2 _03034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_2_3__f_clock_a_I clknet_0_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10855_ _04012_ _05285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_72_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07779__I _02360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13574_ _01453_ clknet_leaf_20_clock u2.mem\[194\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_10786_ _05244_ _01003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12525_ _00404_ clknet_leaf_188_clock u2.mem\[25\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07464__A1 _02933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12588__CLK clknet_leaf_190_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_119_clock_I clknet_5_15_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12456_ _00335_ clknet_leaf_126_clock u2.mem\[20\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07216__A1 _02672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11407_ _05634_ _01234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08264__I0 _03570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12387_ _00266_ clknet_leaf_77_clock u2.mem\[16\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11030__S _05395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07767__A2 _03146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10071__I0 _04801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11338_ _05510_ _05591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12072__D data_in_trans\[11\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11269_ _05504_ _05548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09435__S _04406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13008_ _00887_ clknet_leaf_240_clock u2.mem\[55\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07463__B _02745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09234__I _04170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09516__I0 _04378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10126__I1 u2.mem\[46\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11323__I0 _05554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_1_0_clock_I clknet_4_0_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07500_ u2.mem\[40\]\[7\] _02785_ _02786_ u2.mem\[30\]\[7\] _02972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08480_ _03723_ u2.mem\[8\]\[15\] _03793_ _03797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13363__CLK clknet_leaf_358_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07431_ _02901_ _02902_ _02903_ _02904_ _02905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_91_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07362_ _02581_ _02837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11626__I1 u2.mem\[176\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09101_ _04181_ _04197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_149_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06313_ u2.mem\[189\]\[3\] _01650_ _01652_ u2.mem\[176\]\[3\] _01817_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07293_ u2.mem\[23\]\[3\] _02680_ _02681_ u2.mem\[22\]\[3\] _02769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11004__I _05334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09032_ _04149_ _00344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06244_ u2.mem\[184\]\[1\] _01625_ _01749_ _01750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08514__S _03818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08255__I0 _03561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06175_ _01681_ _01682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07758__A2 _03055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09934_ _04685_ u2.mem\[42\]\[1\] _04719_ _04721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09345__S _04346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09755__I0 _04609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09865_ _04674_ _00652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06718__B1 _02013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11562__I0 _05711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06718__C2 u2.mem\[189\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08816_ _03935_ u2.mem\[16\]\[13\] _04005_ _04007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09796_ _04609_ u2.mem\[38\]\[13\] _04633_ _04635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07391__B1 _02820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09507__I0 _04369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07930__A2 _02559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08747_ _03965_ _00243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08678_ _03922_ _00217_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11865__I1 u2.mem\[191\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07629_ _02443_ _03099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06497__A2 _01917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07694__B2 u2.mem\[30\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07599__I _02581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12730__CLK clknet_leaf_43_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10640_ _05154_ _00947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08238__A3 _03633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06436__C _01934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08494__I0 _03806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_120_clock_I clknet_5_15_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10954__S _05336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10571_ _05111_ _00921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12310_ _00189_ clknet_leaf_99_clock u2.mem\[11\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07997__A2 _03458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13290_ _01169_ clknet_leaf_354_clock u2.mem\[151\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06008__I _01512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12880__CLK clknet_leaf_230_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12241_ _00120_ clknet_leaf_227_clock u2.mem\[7\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08246__I0 _03552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12172_ _00051_ clknet_leaf_210_clock u2.mem\[3\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11785__S _05866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11123_ _05455_ _01129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09746__I0 _04602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11054_ _05411_ _05402_ _05412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_49_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11553__I0 _05717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_254_clock clknet_5_23_0_clock clknet_leaf_254_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_49_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10005_ _04334_ _04760_ _04761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09054__I data_in_trans\[12\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12260__CLK clknet_leaf_70_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13386__CLK clknet_leaf_306_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_45_clock_I clknet_5_6_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11305__I0 _05550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_269_clock clknet_5_22_0_clock clknet_leaf_269_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11956_ _05974_ _01443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10907_ _05318_ _05319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06488__A2 _01970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11887_ u2.mem\[192\]\[4\] _03507_ _05932_ _05935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11608__I1 u2.mem\[175\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10838_ _05273_ _03986_ _05274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_160_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07437__A1 u2.mem\[28\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08485__I0 _03798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12067__D net22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10864__S _05287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10769_ _05200_ u2.mem\[62\]\[2\] _05232_ _05235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13557_ _01436_ clknet_leaf_19_clock u2.mem\[193\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07988__A2 _02627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12508_ _00387_ clknet_leaf_180_clock u2.mem\[24\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13488_ _01367_ clknet_leaf_298_clock u2.mem\[184\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12439_ _00318_ clknet_leaf_127_clock u2.mem\[19\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10663__I _05151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06660__A2 _02125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_207_clock clknet_5_29_0_clock clknet_leaf_207_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_160_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11695__S _05809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06412__A2 _01912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_322_clock_I clknet_5_18_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07980_ u2.mem\[9\]\[15\] _03302_ _03303_ u2.mem\[25\]\[15\] _03444_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12603__CLK clknet_leaf_196_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06931_ _02409_ _02410_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_122_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11494__I _05605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09650_ _04491_ u2.mem\[35\]\[12\] _04537_ _04538_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06862_ col_select_trans\[5\].data_sync _02025_ _02341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_clock clock clknet_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08601_ _03826_ u2.mem\[11\]\[12\] _03872_ _03873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08960__I1 u2.mem\[20\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09581_ _04176_ _04498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06793_ u2.mem\[177\]\[4\] _02091_ _02088_ u2.mem\[193\]\[4\] _02274_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08532_ _03722_ _03833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12753__CLK clknet_leaf_230_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07125__B1 _02603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08463_ _03787_ _00137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06479__A2 _01955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07414_ _02522_ _02888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08394_ _03715_ u2.mem\[6\]\[13\] _03743_ _03745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07345_ _02791_ _02803_ _02812_ _02819_ _02820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_52_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08476__I0 _03715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10774__S _05237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07428__B2 u2.mem\[62\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08244__S _03635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07276_ _02748_ _02749_ _02750_ _02751_ _02752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_148_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09015_ _04135_ _04136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06227_ u2.mem\[193\]\[1\] _01731_ _01732_ u2.mem\[168\]\[1\] _01733_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12133__CLK clknet_leaf_14_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10573__I _05094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06651__A2 _02044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13259__CLK clknet_leaf_311_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06158_ _01564_ _01665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06403__A2 _01681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06089_ _01587_ _01596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09075__S _04182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09917_ _04604_ _04709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11535__I0 _05715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08156__A2 _03583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09848_ _04576_ u2.mem\[40\]\[3\] _04661_ _04665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06167__A1 u2.mem\[144\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06167__B2 u2.mem\[182\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06706__A3 _02189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09779_ _04625_ _00615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11810_ _05768_ _05886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12790_ _00669_ clknet_leaf_71_clock u2.mem\[41\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11741_ _05833_ u2.mem\[183\]\[3\] _05840_ _05844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11672_ _05786_ u2.mem\[179\]\[0\] _05801_ _05802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07122__I _02600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10623_ _05144_ _00940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13411_ _01290_ clknet_leaf_341_clock u2.mem\[172\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08467__I0 _03698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_271_clock_I clknet_5_20_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10684__S _05179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13342_ _01221_ clknet_leaf_4_clock u2.mem\[160\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10554_ _05099_ u2.mem\[57\]\[2\] _05095_ _05100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06642__A2 _02052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13273_ _01152_ clknet_leaf_9_clock u2.mem\[149\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10485_ _05007_ u2.mem\[55\]\[6\] _05056_ _05059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12224_ _00103_ clknet_leaf_231_clock u2.mem\[6\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12626__CLK clknet_leaf_170_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11774__I0 _05837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12155_ _00034_ clknet_leaf_204_clock u2.mem\[2\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08888__I _04050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_2_0_clock clknet_0_clock clknet_3_2_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_116_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_193_clock clknet_5_31_0_clock clknet_leaf_193_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07792__I _02460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11106_ _05420_ u2.mem\[144\]\[0\] _05445_ _05446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12086_ mem_write_n_trans.A clknet_leaf_288_clock mem_write_n_trans.data_sync vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11526__I0 _05707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12776__CLK clknet_leaf_130_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11037_ _05401_ _01097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06201__I _01707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12006__CLK clknet_leaf_312_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11829__I1 u2.mem\[189\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12988_ _00867_ clknet_leaf_257_clock u2.mem\[54\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11939_ _05220_ u2.mem\[193\]\[11\] _05960_ _05964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_131_clock clknet_5_12_0_clock clknet_leaf_131_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08128__I _03545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06330__A1 u2.mem\[154\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07032__I _02510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06330__B2 u2.mem\[162\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12156__CLK clknet_leaf_205_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08458__I0 _03681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07130_ u2.mem\[18\]\[0\] _02606_ _02608_ u2.mem\[19\]\[0\] _02609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_146_clock clknet_5_24_0_clock clknet_leaf_146_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_9_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10393__I _05000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07061_ _02539_ _02540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07830__A1 _03287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06012_ u2.driver_mem\[0\] _01517_ _01519_ _01520_ _01521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_138_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06397__A1 u2.mem\[152\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07594__B1 _02907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07963_ u2.mem\[54\]\[15\] _02509_ _02511_ u2.mem\[55\]\[15\] _03427_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11517__I0 _05674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09702_ _04126_ _04569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06914_ _02378_ _02391_ _02392_ _02393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_68_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07894_ u2.mem\[9\]\[13\] _03302_ _03303_ u2.mem\[25\]\[13\] _03360_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06149__A1 _01561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07346__B1 _02667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09623__S _04522_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07897__A1 u2.mem\[23\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09633_ _04528_ _00566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06845_ u2.mem\[194\]\[5\] _02133_ _02134_ u2.mem\[190\]\[5\] _02325_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10769__S _05232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07897__B2 u2.mem\[22\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11952__I _05971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09564_ _04486_ _00539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06776_ u2.mem\[165\]\[3\] _02075_ _02078_ u2.mem\[163\]\[3\] _02258_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_5_4_0_clock clknet_4_2_0_clock clknet_5_4_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_43_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08515_ _03821_ _00155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09495_ _04442_ _04443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08697__I0 _03935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08446_ _03777_ _03778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_71_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06321__A1 u2.mem\[159\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06321__B2 u2.mem\[149\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08377_ _03735_ _00103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08449__I0 _03664_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06872__A2 _02350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13081__CLK clknet_leaf_40_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07328_ _02794_ _02797_ _02800_ _02802_ _02803_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__12649__CLK clknet_leaf_111_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08074__A1 _01962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11399__I _05507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07259_ _02720_ _02725_ _02730_ _02735_ _02736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__06624__A2 _02037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10009__S _04762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10270_ _04893_ u2.mem\[50\]\[3\] _04923_ _04927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11756__I0 _05833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06388__A1 u2.mem\[145\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06388__B2 u2.mem\[168\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_218_clock_I clknet_5_28_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12029__CLK clknet_2_2__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11133__A1 _05295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07117__I _02595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12911_ _00790_ clknet_leaf_157_clock u2.mem\[49\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10679__S _05174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07888__B2 u2.mem\[62\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12842_ _00721_ clknet_leaf_139_clock u2.mem\[44\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12773_ _00652_ clknet_leaf_79_clock u2.mem\[40\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13424__CLK clknet_leaf_347_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11724_ _03670_ _05833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06312__A1 u2.mem\[174\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06312__B2 u2.mem\[150\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11655_ _05667_ _05790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_63_clock clknet_5_9_0_clock clknet_leaf_63_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06863__A2 _02024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07787__I _02427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10247__I0 _04911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11303__S _05568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10606_ _05101_ u2.mem\[58\]\[3\] _05131_ _05135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11586_ _05662_ _05746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13574__CLK clknet_leaf_20_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10798__I1 u2.mem\[62\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13325_ _01204_ clknet_leaf_342_clock u2.mem\[157\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06615__A2 _02053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10537_ _05020_ u2.mem\[56\]\[12\] _05088_ _05089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08860__I0 _04037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_78_clock clknet_5_8_0_clock clknet_leaf_78_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_48_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09708__S _04567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13256_ _01135_ clknet_leaf_311_clock u2.mem\[146\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10468_ _05027_ u2.mem\[54\]\[15\] _05045_ _05049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12207_ _00086_ clknet_leaf_229_clock u2.mem\[5\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10941__I _05339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13187_ _01066_ clknet_leaf_274_clock u2.mem\[134\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06379__A1 u2.mem\[180\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10399_ _05005_ u2.mem\[53\]\[5\] _05002_ _05006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07576__B1 _02891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06379__B2 u2.mem\[150\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12138_ _01464_ clknet_leaf_38_clock u2.driver_mem\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07040__A2 _02403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11973__S _05980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12080__D data_in_trans\[15\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12069_ net8 clknet_2_0__leaf_clock_a data_in_trans\[10\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07879__B2 u2.mem\[36\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06630_ _02114_ _02115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_16_clock clknet_5_2_0_clock clknet_leaf_16_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_20_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06561_ _02032_ _02036_ _02046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10388__I _04134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08300_ _03675_ _03676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09280_ _04285_ u2.mem\[26\]\[15\] _04305_ _04309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06303__A1 _01769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06492_ _01976_ _01970_ _01977_ _01978_ _01463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08231_ _03579_ u2.mem\[3\]\[15\] _03624_ _03628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10238__I0 _04904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08162_ _03550_ u2.mem\[2\]\[2\] _03585_ _03588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08056__A1 _03511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_167_clock_I clknet_5_26_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07113_ _02418_ _02420_ _02404_ _02547_ _02592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_88_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08093_ u2.driver_enable output_active_hold\[1\] output_active_hold\[0\] _03538_
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06606__A2 _02015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12941__CLK clknet_leaf_256_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11012__I _05342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07044_ _02522_ _02523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08603__I0 _03829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11363__A1 _03487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07567__B1 _02882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08321__I _03692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08995_ _04118_ _04119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11883__S _05932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07582__A3 _03045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07946_ u2.mem\[39\]\[14\] _03321_ _03322_ u2.mem\[48\]\[14\] _03411_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_5_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06790__A1 _02245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input27_I mem_address_a[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07877_ u2.mem\[54\]\[13\] _02509_ _02511_ u2.mem\[55\]\[13\] _03343_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10499__S _05066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_27_0_clock clknet_4_13_0_clock clknet_5_27_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_110_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12321__CLK clknet_leaf_158_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10713__I1 u2.mem\[61\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13447__CLK clknet_leaf_343_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09616_ _04518_ _00559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06828_ u2.mem\[184\]\[5\] _02072_ _01994_ _02308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09547_ _04473_ u2.mem\[33\]\[4\] _04474_ _04475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06759_ u2.mem\[187\]\[3\] _02186_ _02187_ u2.mem\[192\]\[3\] _02241_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_70_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09478_ _04380_ u2.mem\[31\]\[10\] _04429_ _04432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08429_ _03702_ u2.mem\[7\]\[10\] _03764_ _03767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06845__A2 _02133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06725__B _01995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11440_ _04120_ _05645_ _05654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_36_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08047__A1 _01809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09095__I0 _04158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11371_ _05591_ u2.mem\[160\]\[3\] _05608_ _05612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_1497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10322_ _04956_ _00827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13110_ _00989_ clknet_leaf_19_clock u2.mem\[61\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07270__A2 _02480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13041_ _00920_ clknet_leaf_321_clock u2.mem\[57\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09398__I1 u2.mem\[29\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10253_ _04608_ _04916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07022__A2 _02495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10184_ _04871_ _00774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06781__A1 u2.mem\[150\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06781__B2 u2.mem\[174\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07730__B1 _03092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12814__CLK clknet_leaf_220_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12825_ _00704_ clknet_leaf_136_clock u2.mem\[43\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10468__I0 _05027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08607__S _03872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12756_ _00635_ clknet_leaf_69_clock u2.mem\[39\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11707_ _05794_ u2.mem\[181\]\[3\] _05818_ _05822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06836__A2 _02103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12687_ _00566_ clknet_leaf_175_clock u2.mem\[35\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12964__CLK clknet_leaf_109_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08038__A1 _03497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09086__I0 _04145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08406__I _03753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11638_ _05746_ u2.mem\[177\]\[0\] _05779_ _05780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07310__I _02405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12075__D net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11569_ _05736_ _01294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13308_ _01187_ clknet_leaf_353_clock u2.mem\[154\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07261__A2 _02633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13239_ _01118_ clknet_leaf_284_clock u2.mem\[143\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09237__I _04173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08141__I _03545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07800_ _02479_ _03267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08780_ mem_address_trans\[4\].data_sync _03984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_38_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06772__A1 u2.mem\[184\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09173__S _04236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07731_ u2.mem\[6\]\[10\] _03094_ _03095_ u2.mem\[47\]\[10\] _03200_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_66_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07316__A3 _02787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_93_clock_I clknet_5_10_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10112__S _04825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07662_ _02558_ _03132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12494__CLK clknet_leaf_181_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07721__B1 _03073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09401_ _04357_ _04385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_4_1492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06613_ _02007_ _02080_ _02098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07593_ _03054_ _03057_ _03060_ _03063_ _03064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_59_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09313__I1 u2.mem\[27\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10459__I0 _05018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09332_ _04340_ _00453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06544_ _02023_ _02028_ _02029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08517__S _03818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11120__I1 u2.mem\[145\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09263_ _04299_ _00425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06475_ _01962_ _01955_ _01963_ _01965_ _01459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08214_ _03618_ _00057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09194_ _04253_ _00402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09077__I0 _04128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08316__I _03688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08145_ _03575_ u2.mem\[1\]\[13\] _03573_ _03576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10631__I0 _05126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07252__A2 _02606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08076_ _03525_ _03519_ _03526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_162_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07027_ u2.mem\[50\]\[0\] _02503_ _02505_ u2.mem\[51\]\[0\] _02506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06460__B1 _01952_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11187__I1 u2.mem\[149\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08051__I _03493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07095__C _02568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08978_ _04035_ u2.mem\[20\]\[9\] _04107_ _04109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06763__A1 u2.mem\[154\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06763__B2 u2.mem\[162\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09001__I0 _04119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07929_ _03378_ _03383_ _03388_ _03393_ _03394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_99_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10022__S _04767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10940_ _04126_ _05339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06439__C _01934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10871_ _03582_ _05295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_77_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_1_0_clock clknet_3_0_0_clock clknet_4_1_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_164_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12987__CLK clknet_leaf_248_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09304__I1 u2.mem\[27\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12610_ _00489_ clknet_leaf_173_clock u2.mem\[30\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12541_ _00420_ clknet_leaf_188_clock u2.mem\[26\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12217__CLK clknet_leaf_53_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12472_ _00351_ clknet_leaf_121_clock u2.mem\[21\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07491__A2 _02920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11788__S _05866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11423_ _05635_ u2.mem\[163\]\[5\] _05637_ _05644_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09258__S _04295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10622__I0 _05117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11354_ _05601_ _01214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08162__S _03585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07243__A2 _02717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12367__CLK clknet_leaf_223_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10305_ _04891_ u2.mem\[51\]\[2\] _04944_ _04947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11285_ _05558_ _05559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_140_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10236_ _04591_ _04904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_1565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13024_ _00903_ clknet_leaf_246_clock u2.mem\[56\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10167_ _04817_ u2.mem\[47\]\[15\] _04856_ _04860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09791__I1 u2.mem\[38\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06754__A1 u2.mem\[169\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_115_clock_I clknet_5_14_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06754__B2 u2.mem\[147\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06410__S _01510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10098_ _04821_ _00738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11028__S _05395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_1_0_clock_I clknet_3_0_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07703__B1 _03115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07305__I _02360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12808_ _00687_ clknet_leaf_139_clock u2.mem\[42\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12739_ _00618_ clknet_leaf_65_clock u2.mem\[38\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06260_ _01759_ _01760_ _01765_ _01766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_148_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13142__CLK clknet_leaf_23_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06191_ _01567_ _01665_ _01678_ _01698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_117_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10613__I0 _05108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07234__A2 _02657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09950_ _04700_ u2.mem\[42\]\[8\] _04729_ _04730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13292__CLK clknet_leaf_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11169__I1 u2.mem\[148\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08901_ _04063_ _00299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08800__S _03995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09881_ _04684_ _00658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08832_ _04018_ _00275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06745__A1 u2.mem\[153\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06745__B2 u2.mem\[160\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08763_ _03974_ _00250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07714_ u2.mem\[60\]\[10\] _03055_ _03056_ u2.mem\[62\]\[10\] _03183_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08694_ _03932_ u2.mem\[13\]\[12\] _03933_ _03934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07645_ _02510_ _03115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07576_ u2.mem\[14\]\[8\] _02890_ _02891_ u2.mem\[12\]\[8\] _03047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_317_clock_I clknet_5_18_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09315_ _04281_ u2.mem\[27\]\[13\] _04328_ _04330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06527_ _02011_ _02001_ _02012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10576__I _03696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09246_ _04289_ _04290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06458_ u2.mem\[194\]\[7\] _01946_ _01952_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09177_ _04225_ _04241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06389_ u2.mem\[187\]\[5\] _01632_ _01635_ u2.mem\[192\]\[5\] _01891_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08128_ _03545_ _03564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10604__I0 _05099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07225__A2 _02475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08273__I1 u2.mem\[4\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08059_ _03513_ _03508_ _03514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06984__A1 _02440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09806__S _04639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11070_ _05421_ _05422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09222__I0 _04272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10021_ _04770_ _00712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06736__B2 u2.mem\[161\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11580__I1 u2.mem\[173\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13015__CLK clknet_leaf_323_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09525__I1 u2.mem\[32\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11972_ _05983_ _01450_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10923_ _05328_ _01056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10854_ _05284_ _01031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13165__CLK clknet_leaf_264_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11096__I0 _05428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13573_ _01452_ clknet_leaf_20_clock u2.mem\[194\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10785_ _05216_ u2.mem\[62\]\[9\] _05242_ _05244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11796__A1 _04310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12524_ _00403_ clknet_leaf_187_clock u2.mem\[25\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10843__I0 _05194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07464__A2 _02934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12455_ _00334_ clknet_leaf_127_clock u2.mem\[20\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_41_clock_I clknet_5_6_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07795__I _02470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11311__S _05567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11406_ _05633_ u2.mem\[162\]\[4\] _05624_ _05634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07216__A2 _02679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12386_ _00265_ clknet_leaf_224_clock u2.mem\[16\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08264__I1 u2.mem\[4\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11337_ _05590_ _01208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11268_ _05547_ _01182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07519__A3 _02985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13007_ _00886_ clknet_leaf_240_clock u2.mem\[55\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10219_ _04892_ _00788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07744__B _03211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11199_ _05500_ u2.mem\[150\]\[0\] _05502_ _05503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06727__A1 u2.mem\[150\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07924__B1 _02523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_266_clock_I clknet_5_23_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09516__I1 u2.mem\[32\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11323__I1 u2.mem\[157\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13508__CLK clknet_leaf_331_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07430_ u2.mem\[57\]\[5\] _02828_ _02829_ u2.mem\[41\]\[5\] _02904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_5_0_clock_I clknet_4_2_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07361_ _02579_ _02836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12532__CLK clknet_leaf_98_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09100_ _04196_ _00365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06312_ u2.mem\[174\]\[3\] _01656_ _01666_ u2.mem\[150\]\[3\] _01660_ u2.mem\[181\]\[3\]
+ _01816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_07292_ _02764_ _02765_ _02766_ _02767_ _02768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_143_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07455__A2 _02866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09031_ _04148_ u2.mem\[21\]\[6\] _04141_ _04149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06243_ _01553_ _01749_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07207__A2 _02606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06174_ _01581_ _01599_ _01681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12682__CLK clknet_leaf_127_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09933_ _04720_ _00674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13038__CLK clknet_leaf_248_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09864_ _04599_ u2.mem\[40\]\[10\] _04671_ _04674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06718__A1 u2.mem\[176\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09425__I _04395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06718__B2 u2.mem\[172\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11562__I1 u2.mem\[172\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08815_ _04006_ _00270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09795_ _04634_ _00622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07391__A1 _01843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09507__I1 u2.mem\[32\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08746_ _03908_ u2.mem\[15\]\[1\] _03963_ _03965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12062__CLK clknet_leaf_302_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13188__CLK clknet_leaf_270_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08677_ _03921_ u2.mem\[13\]\[7\] _03915_ _03922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08191__I0 _03579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07628_ _01954_ _03013_ _03053_ _03098_ _01500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06351__C1 u2.mem\[165\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07559_ u2.mem\[1\]\[8\] _03028_ _03029_ u2.mem\[7\]\[8\] _03030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_41_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10570_ _05110_ u2.mem\[57\]\[7\] _05104_ _05111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09229_ _04277_ _00413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12240_ _00119_ clknet_leaf_227_clock u2.mem\[7\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06406__B1 _01679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12171_ _00050_ clknet_leaf_209_clock u2.mem\[3\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11950__A1 _03582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11122_ _05424_ u2.mem\[145\]\[1\] _05453_ _05455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08440__S _03769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11053_ _03903_ _05411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_67_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07564__B _02978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06959__I _02370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06709__A1 u2.mem\[180\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06709__B2 u2.mem\[150\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10004_ _04440_ _04760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11553__I1 u2.mem\[171\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09271__S _04300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11305__I1 u2.mem\[156\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11955_ _05907_ u2.mem\[194\]\[1\] _05972_ _05974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07134__A1 _02466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08182__I0 _03570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10906_ _04095_ _05317_ _05318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07685__A2 _03153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11886_ _05934_ _01413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06627__C _02111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10837_ mem_address_trans\[6\].data_sync _05273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13556_ _01435_ clknet_leaf_18_clock u2.mem\[193\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08615__S _03880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10768_ _05234_ _00995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12507_ _00386_ clknet_leaf_179_clock u2.mem\[24\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10944__I _04130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13487_ _01366_ clknet_leaf_296_clock u2.mem\[184\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11041__S _05404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10699_ _05119_ u2.mem\[60\]\[11\] _05184_ _05188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12438_ _00317_ clknet_leaf_87_clock u2.mem\[19\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11976__S _05985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10880__S _05297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12369_ _00248_ clknet_leaf_223_clock u2.mem\[15\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_361_clock clknet_5_0_0_clock clknet_leaf_361_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06930_ _02352_ _02376_ _02409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_132_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12085__CLK clknet_2_2__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I col_select_a[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13330__CLK clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06861_ row_select_trans\[0\].data_sync row_select_trans\[2\].data_sync _02340_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06176__A2 _01641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08600_ _03856_ _03872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09580_ _04497_ _00544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06792_ u2.mem\[151\]\[4\] _02084_ _02086_ u2.mem\[158\]\[4\] u2.mem\[168\]\[4\]
+ _02093_ _02273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_83_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08531_ _03832_ _00160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07125__A1 u2.mem\[52\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08173__I0 _03561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13480__CLK clknet_leaf_289_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08462_ _03689_ u2.mem\[8\]\[7\] _03783_ _03787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07413_ _02520_ _02887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08393_ _03744_ _00110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11015__I _05345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07344_ _02813_ _02814_ _02815_ _02818_ _02819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_10_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06109__I _01580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08476__I1 u2.mem\[8\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07275_ u2.mem\[58\]\[3\] _02495_ _02500_ u2.mem\[36\]\[3\] _02751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09014_ _04134_ _04135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06226_ _01589_ _01732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_314_clock clknet_5_19_0_clock clknet_leaf_314_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_128_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_0_0_clock clknet_4_0_0_clock clknet_5_0_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_06157_ _01663_ _01664_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12428__CLK clknet_leaf_180_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07600__A2 _03069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08260__S _03645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06088_ _01594_ _01595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_329_clock clknet_5_7_0_clock clknet_leaf_329_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09916_ _04708_ _00669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11535__I1 u2.mem\[170\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09847_ _04664_ _00644_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_9_clock_I clknet_5_1_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08994__I _04117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09778_ _04583_ u2.mem\[38\]\[5\] _04623_ _04625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08729_ _03928_ u2.mem\[14\]\[10\] _03952_ _03955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08164__I0 _03552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11126__S _05453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11740_ _05843_ _01358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11671_ _05800_ _05801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10965__S _05356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_214_clock_I clknet_5_28_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13410_ _01289_ clknet_leaf_305_clock u2.mem\[171\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10622_ _05117_ u2.mem\[58\]\[10\] _05141_ _05144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08467__I1 u2.mem\[8\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13341_ _01220_ clknet_leaf_3_clock u2.mem\[160\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10764__I _05231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10553_ _04994_ _05099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13203__CLK clknet_leaf_280_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13272_ _01151_ clknet_5_0_0_clock u2.mem\[148\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10484_ _05058_ _00887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12223_ _00102_ clknet_leaf_231_clock u2.mem\[6\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11774__I1 u2.mem\[185\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12154_ _00033_ clknet_leaf_56_clock u2.mem\[1\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13353__CLK clknet_leaf_358_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11105_ _05444_ _05445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_68_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10205__S _04880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12085_ net34 clknet_2_2__leaf_clock_a mem_write_n_trans.A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11526__I1 u2.mem\[170\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11036_ _05392_ u2.mem\[139\]\[5\] _05394_ _05401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07355__B2 u2.mem\[41\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10004__I _04440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12987_ _00866_ clknet_leaf_248_clock u2.mem\[54\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11036__S _05394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07658__A2 _03126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11938_ _05963_ _01436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07313__I _02427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12078__D data_in_trans\[14\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11869_ _05913_ u2.mem\[191\]\[4\] _05917_ _05923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06330__A2 _01698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11462__I0 _05668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10674__I _05173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13539_ _01418_ clknet_leaf_34_clock u2.mem\[192\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06094__A1 _01599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07060_ _02455_ _02537_ _02538_ _02484_ _02539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__07291__B1 _02587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08144__I _03531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07830__A2 _03290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06011_ _01503_ _01520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06397__A2 _01712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10115__S _04830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07962_ u2.mem\[50\]\[15\] _02503_ _02505_ u2.mem\[51\]\[15\] _03426_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12720__CLK clknet_leaf_236_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_13_0_clock_I clknet_4_6_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09701_ _04568_ _00594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06913_ _02348_ _02350_ _02392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_136_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07893_ u2.mem\[29\]\[13\] _03299_ _03300_ u2.mem\[11\]\[13\] _03359_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07346__A1 u2.mem\[61\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08394__I0 _03715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_163_clock_I clknet_5_26_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09632_ _04473_ u2.mem\[35\]\[4\] _04527_ _04528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06844_ u2.mem\[144\]\[5\] _02114_ _02116_ u2.mem\[182\]\[5\] _02324_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07897__A2 _02596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12870__CLK clknet_leaf_83_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09563_ _04485_ u2.mem\[33\]\[9\] _04483_ _04486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06775_ u2.mem\[151\]\[3\] _02084_ _02086_ u2.mem\[158\]\[3\] u2.mem\[193\]\[3\]
+ _02088_ _02257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_167_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08514_ _03820_ u2.mem\[9\]\[9\] _03818_ _03821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09494_ _03983_ _04441_ _04442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_110_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08319__I data_in_trans\[8\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08445_ _03630_ _03542_ _03776_ _03777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_24_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10785__S _05242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13226__CLK clknet_leaf_279_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08376_ _03681_ u2.mem\[6\]\[5\] _03733_ _03735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07327_ u2.mem\[3\]\[4\] _02801_ _02745_ _02802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_253_clock clknet_5_22_0_clock clknet_leaf_253_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_143_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08074__A2 _03517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12250__CLK clknet_leaf_57_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08054__I data_in_trans\[5\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_23_0_clock clknet_4_11_0_clock clknet_5_23_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07258_ _02731_ _02732_ _02733_ _02734_ _02735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_clkbuf_leaf_88_clock_I clknet_5_10_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06209_ u2.mem\[152\]\[0\] _01713_ _01715_ u2.mem\[148\]\[0\] _01716_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07189_ _02560_ _02667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_151_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11756__I1 u2.mem\[184\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_268_clock clknet_5_22_0_clock clknet_leaf_268_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_160_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10025__S _04772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07337__A1 _02804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08385__I0 _03698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11133__A2 _05443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12910_ _00789_ clknet_leaf_202_clock u2.mem\[49\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10192__I0 _04801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12841_ _00720_ clknet_leaf_138_clock u2.mem\[44\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_206_clock clknet_5_29_0_clock clknet_leaf_206_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12772_ _00651_ clknet_leaf_91_clock u2.mem\[40\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07133__I _02611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11723_ _05832_ _01352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10695__S _05184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06312__A2 _01656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06972__I _02407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11654_ _05789_ _01326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11444__I0 _05627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10605_ _05134_ _00932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11585_ _05745_ _01301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06076__A1 _01582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13324_ _01203_ clknet_leaf_342_clock u2.mem\[157\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07273__B1 _02649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10536_ _05072_ _05088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07812__A2 _03120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13255_ _01134_ clknet_leaf_295_clock u2.mem\[146\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12743__CLK clknet_leaf_53_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10467_ _05048_ _00880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12206_ _00085_ clknet_leaf_212_clock u2.mem\[5\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13186_ _01065_ clknet_leaf_276_clock u2.mem\[134\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_1506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07576__A1 u2.mem\[14\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10398_ _05004_ _05005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07576__B2 u2.mem\[12\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12137_ _01463_ clknet_leaf_38_clock u2.driver_mem\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07040__A3 _02383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07308__I _02395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12893__CLK clknet_leaf_214_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12068_ data_in_trans\[9\].A clknet_leaf_33_clock data_in_trans\[9\].data_sync vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08376__I0 _03681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11019_ _05390_ u2.mem\[138\]\[4\] _05381_ _05391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10183__I0 _04792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12123__CLK clknet_leaf_37_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13249__CLK clknet_leaf_285_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06560_ _02044_ _02045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10635__A1 _04311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06491_ u2.mem\[193\]\[14\] _01917_ _01919_ u2.mem\[192\]\[14\] _01920_ _01978_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08230_ _03627_ _00064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12273__CLK clknet_leaf_165_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06882__I _02360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08161_ _03587_ _00035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07112_ _02590_ _02591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07264__B1 _02436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08092_ output_active_hold\[3\] output_active_hold\[2\] _03537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07803__A2 _03111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07043_ _02429_ _02445_ _02446_ _02493_ _02522_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_118_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08603__I1 u2.mem\[11\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09800__I0 _04615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11363__A2 _05606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08994_ _04117_ _04118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06775__C1 u2.mem\[193\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09634__S _04527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07582__A4 _03052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07945_ u2.mem\[5\]\[14\] _02627_ _02629_ u2.mem\[38\]\[14\] _03410_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08367__I0 _03664_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06790__A2 _02249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10174__I0 _04782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07876_ u2.mem\[50\]\[13\] _02503_ _02505_ u2.mem\[51\]\[13\] _03342_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09615_ _04494_ u2.mem\[34\]\[13\] _04516_ _04518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06827_ u2.mem\[167\]\[5\] _02060_ _02062_ u2.mem\[183\]\[5\] _02307_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10579__I _03700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08119__I0 _03557_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09546_ _04464_ _04474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_37_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08049__I data_in_trans\[4\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06758_ u2.mem\[159\]\[3\] _02174_ _02176_ u2.mem\[149\]\[3\] _02240_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12616__CLK clknet_leaf_113_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11674__I0 _05790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09477_ _04431_ _00507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06689_ u2.mem\[145\]\[1\] _02082_ _02094_ u2.mem\[168\]\[1\] _02173_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08428_ _03766_ _00123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_192_clock clknet_5_31_0_clock clknet_leaf_192_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09619__I0 _04498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08359_ _03723_ u2.mem\[5\]\[15\] _03711_ _03724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12766__CLK clknet_leaf_203_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07255__B1 _02619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11370_ _05611_ _01220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08713__S _03942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10321_ _04907_ u2.mem\[51\]\[9\] _04954_ _04956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13040_ _00919_ clknet_leaf_320_clock u2.mem\[57\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10252_ _04915_ _00798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10183_ _04792_ u2.mem\[48\]\[4\] _04870_ _04871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_130_clock clknet_5_14_0_clock clknet_leaf_130_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_117_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06781__A2 _02047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_1_0_clock_I clknet_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10165__I0 _04815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06967__I _02432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11901__I1 _03523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_145_clock clknet_5_24_0_clock clknet_leaf_145_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10489__I _05050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07730__B2 u2.mem\[4\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12824_ _00703_ clknet_leaf_137_clock u2.mem\[43\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12296__CLK clknet_leaf_120_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13541__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11665__I0 _05796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12755_ _00634_ clknet_leaf_64_clock u2.mem\[39\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08530__I0 _03831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06916__B _02393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07798__I _02476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06297__A1 u2.mem\[191\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11706_ _05821_ _01346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06297__B2 u2.mem\[179\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12686_ _00565_ clknet_leaf_193_clock u2.mem\[35\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11417__I0 _05629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11637_ _05778_ _05779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_leaf_111_clock_I clknet_5_14_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07246__B1 _02582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11568_ _05717_ u2.mem\[172\]\[4\] _05730_ _05736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13307_ _01186_ clknet_leaf_359_clock u2.mem\[154\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10952__I _04138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10519_ _05001_ u2.mem\[56\]\[4\] _05078_ _05079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11499_ _05668_ u2.mem\[168\]\[1\] _05692_ _05694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13238_ _01117_ clknet_leaf_284_clock u2.mem\[143\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07549__B2 u2.mem\[30\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11984__S _05971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12091__D net23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13169_ _01048_ clknet_leaf_265_clock u2.mem\[131\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07038__I _02516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08349__I0 _03715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13071__CLK clknet_leaf_240_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07730_ u2.mem\[8\]\[10\] _03091_ _03092_ u2.mem\[4\]\[10\] _03199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10156__I0 _04806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_36_clock_I clknet_5_4_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10856__A1 _05285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07661_ _03105_ _03110_ _03119_ _03130_ _03131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_26_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07721__A1 u2.mem\[28\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07721__B2 u2.mem\[31\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09400_ _04166_ _04384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06612_ _02096_ _02097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07592_ u2.mem\[57\]\[8\] _03061_ _03062_ u2.mem\[41\]\[8\] _03063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09331_ _04258_ u2.mem\[28\]\[3\] _04336_ _04340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11656__I0 _05790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06543_ _02026_ _02027_ _02028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12789__CLK clknet_leaf_71_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06288__A1 _01789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09262_ _04267_ u2.mem\[26\]\[7\] _04295_ _04299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06474_ u2.mem\[193\]\[10\] _01960_ _01948_ u2.mem\[192\]\[10\] _01964_ _01965_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08213_ _03561_ u2.mem\[3\]\[7\] _03614_ _03618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09193_ _04246_ u2.mem\[25\]\[0\] _04252_ _04253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09629__S _04522_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12019__CLK clknet_2_2__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08144_ _03531_ _03575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08075_ data_in_trans\[11\].data_sync _03525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07026_ _02504_ _02505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06460__A1 _01951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08332__I _03701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11894__S _05937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13414__CLK clknet_leaf_342_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_313_clock_I clknet_5_19_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10395__I0 _05001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06212__A1 _01612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08977_ _04108_ _00330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_62_clock clknet_5_9_0_clock clknet_leaf_62_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_25_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07928_ _03389_ _03390_ _03391_ _03392_ _03393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_99_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10303__S _04944_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10147__I0 _04797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07859_ u2.mem\[8\]\[12\] _03324_ _03325_ u2.mem\[4\]\[12\] _03326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07712__A1 _03165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10870_ _04986_ _05294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_77_clock clknet_5_8_0_clock clknet_leaf_77_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_09529_ _04391_ u2.mem\[32\]\[15\] _04458_ _04462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_12540_ _00419_ clknet_leaf_189_clock u2.mem\[26\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07476__B1 _02900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12471_ _00350_ clknet_leaf_122_clock u2.mem\[21\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10973__S _05355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07228__B1 _02646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11422_ _05643_ _01240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11024__A1 _04311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10622__I1 u2.mem\[58\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11353_ _05589_ u2.mem\[159\]\[2\] _05598_ _05601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_15_clock clknet_5_2_0_clock clknet_leaf_15_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10304_ _04946_ _00819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11284_ _04310_ _05527_ _05558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_152_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13023_ _00902_ clknet_leaf_249_clock u2.mem\[56\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13094__CLK clknet_leaf_23_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10235_ _04903_ _00793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10386__I0 _04995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09274__S _04305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10166_ _04859_ _00768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07951__A1 _01976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06754__A2 _02141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11309__S _05567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10138__I0 _04788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10097_ _04782_ u2.mem\[46\]\[0\] _04820_ _04821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07703__B2 u2.mem\[55\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12931__CLK clknet_leaf_232_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_5_0_clock_I clknet_3_2_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12807_ _00686_ clknet_leaf_140_clock u2.mem\[42\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11638__I0 _05746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10999_ _05377_ _01083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12738_ _00617_ clknet_leaf_234_clock u2.mem\[38\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06809__A3 _02288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10310__I0 _04895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07321__I _02470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12086__D mem_write_n_trans.A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10883__S _05297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12669_ _00548_ clknet_leaf_193_clock u2.mem\[34\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_262_clock_I clknet_5_23_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06190_ u2.mem\[147\]\[0\] _01676_ _01680_ u2.mem\[169\]\[0\] _01696_ _01697_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_116_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11778__I _05865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12311__CLK clknet_leaf_118_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10613__I1 u2.mem\[58\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13437__CLK clknet_leaf_350_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06442__A1 u2.mem\[194\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08900_ _04035_ u2.mem\[18\]\[9\] _04061_ _04063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09880_ _04681_ u2.mem\[41\]\[0\] _04683_ _04684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12461__CLK clknet_leaf_196_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08831_ _04017_ u2.mem\[17\]\[1\] _04015_ _04018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07942__A1 u2.mem\[52\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11219__S _05501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08762_ _03923_ u2.mem\[15\]\[8\] _03973_ _03974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07713_ u2.mem\[61\]\[10\] _03132_ _03133_ u2.mem\[63\]\[10\] _03182_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08693_ _03905_ _03933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_113_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11018__I _05348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07644_ _02508_ _03114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10857__I _05286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07575_ u2.mem\[44\]\[8\] _02887_ _02888_ u2.mem\[42\]\[8\] _03046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09314_ _04329_ _00446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06526_ _02009_ _02010_ _02011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08327__I _03697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10301__I0 _04885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11889__S _05932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09245_ _04288_ _04250_ _04289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_107_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06457_ u2.mem\[0\]\[7\] _01951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_21_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06130__C2 u2.mem\[192\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06681__A1 u2.mem\[144\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09176_ _04240_ _00397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06681__B2 u2.mem\[182\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06388_ u2.mem\[145\]\[5\] _01640_ _01732_ u2.mem\[168\]\[5\] _01890_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08127_ _03518_ _03563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10592__I _03717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10604__I1 u2.mem\[58\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06433__A1 u2.mem\[192\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08058_ data_in_trans\[6\].data_sync _03513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06984__A2 _02401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07009_ _02487_ _02445_ _02446_ _02404_ _02488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__09222__I1 u2.mem\[25\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10368__I0 _04916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08997__I _04120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10020_ _04696_ u2.mem\[44\]\[6\] _04767_ _04770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07933__A1 u2.mem\[57\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12954__CLK clknet_leaf_324_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08011__B _01549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09822__S _04649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11971_ _05213_ u2.mem\[194\]\[8\] _05980_ _05983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10922_ _05294_ u2.mem\[133\]\[0\] _05327_ _05328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08438__S _03769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10853_ _05207_ u2.mem\[128\]\[5\] _05277_ _05284_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_13572_ _01451_ clknet_leaf_20_clock u2.mem\[194\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10784_ _05243_ _01002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12523_ _00402_ clknet_leaf_183_clock u2.mem\[25\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11796__A2 _05847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12334__CLK clknet_leaf_206_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06121__B1 _01614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09269__S _04300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06672__A1 _02125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12454_ _00333_ clknet_leaf_85_clock u2.mem\[20\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06980__I _02419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11405_ _05513_ _05633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12385_ _00264_ clknet_leaf_223_clock u2.mem\[16\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07216__A3 _02686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09068__I _04176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06424__A1 u2.mem\[194\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12484__CLK clknet_leaf_105_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11336_ _05589_ u2.mem\[158\]\[2\] _05585_ _05590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10359__I0 _04907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11267_ _05544_ u2.mem\[154\]\[0\] _05546_ _05547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13006_ _00885_ clknet_leaf_259_clock u2.mem\[55\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10218_ _04891_ u2.mem\[49\]\[2\] _04887_ _04892_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07519__A4 _02990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11198_ _05501_ _05502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_leaf_209_clock_I clknet_5_29_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10149_ _04799_ u2.mem\[47\]\[7\] _04846_ _04850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07688__B1 _03095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09531__I _04118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_0 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06360__B1 _01705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11236__A1 _04223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07360_ u2.mem\[29\]\[4\] _02833_ _02834_ u2.mem\[11\]\[4\] _02835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_16_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08147__I _03533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08101__A1 _03483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06311_ u2.mem\[155\]\[3\] _01659_ _01815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07291_ u2.mem\[28\]\[3\] _02585_ _02587_ u2.mem\[31\]\[3\] _02767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_91_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09030_ _04147_ _04148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_5_9_0_clock_I clknet_4_4_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06242_ u2.mem\[171\]\[1\] _01610_ _01614_ u2.mem\[157\]\[1\] _01748_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12827__CLK clknet_leaf_221_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06173_ _01679_ _01680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07000__B _02434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08811__S _04000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09932_ _04681_ u2.mem\[42\]\[0\] _04719_ _04720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09706__I _04130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09863_ _04673_ _00651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07915__A1 u2.mem\[1\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08814_ _03932_ u2.mem\[16\]\[12\] _04005_ _04006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09794_ _04605_ u2.mem\[38\]\[12\] _04633_ _04634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08745_ _03964_ _00242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07679__B1 _03078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08676_ _03688_ _03921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08258__S _03645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07627_ _03064_ _03075_ _03086_ _03097_ _03098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_81_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12357__CLK clknet_leaf_80_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06351__C2 _01645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07558_ _02470_ _03029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06509_ _01993_ _01994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07489_ u2.mem\[18\]\[6\] _02850_ _02851_ u2.mem\[19\]\[6\] _02962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09840__A1 _04224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09228_ _04276_ u2.mem\[25\]\[11\] _04270_ _04277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_5_clock_I clknet_5_0_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_158_clock_I clknet_5_26_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09159_ _04225_ _04231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_107_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06406__A1 u2.mem\[147\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07603__B1 _03073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12170_ _00049_ clknet_leaf_109_clock u2.mem\[2\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06305__I _01808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11121_ _05454_ _01128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11950__A2 _05926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11052_ _05410_ _01103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_210_clock_I clknet_5_29_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10003_ _04759_ _00705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10761__I0 _05229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13132__CLK clknet_leaf_267_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09659__A1 _04095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_18_0_clock clknet_4_9_0_clock clknet_5_18_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_3742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06975__I _02362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11954_ _05973_ _01442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09351__I _04335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07134__A2 _02467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08182__I1 u2.mem\[2\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10905_ _05275_ _05317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_44_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11885_ u2.mem\[192\]\[3\] _03503_ _05932_ _05934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13282__CLK clknet_leaf_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06893__A1 _02339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10836_ _05272_ _01025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13555_ _01434_ clknet_leaf_18_clock u2.mem\[193\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10767_ _05198_ u2.mem\[62\]\[1\] _05232_ _05234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12506_ _00385_ clknet_leaf_121_clock u2.mem\[23\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06645__A1 _02108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07842__B1 _03147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13486_ _01365_ clknet_leaf_298_clock u2.mem\[184\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10698_ _05187_ _00972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12437_ _00316_ clknet_leaf_88_clock u2.mem\[19\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06215__I _01721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08631__S _03890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12368_ _00247_ clknet_leaf_222_clock u2.mem\[15\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11319_ _05550_ u2.mem\[157\]\[2\] _05576_ _05579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12299_ _00178_ clknet_leaf_170_clock u2.mem\[11\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06860_ _02025_ _01989_ _02339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10752__I0 _05222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09462__S _04419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06791_ _01809_ _01995_ _02244_ _02272_ _01477_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08530_ _03831_ u2.mem\[9\]\[14\] _03827_ _03832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06885__I _02363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07125__A2 _02601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08461_ _03786_ _00136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07412_ _02880_ _02883_ _02884_ _02885_ _02886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10200__I _04864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08392_ _03710_ u2.mem\[6\]\[12\] _03743_ _03744_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07343_ u2.mem\[43\]\[4\] _02816_ _02817_ u2.mem\[20\]\[4\] _02818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07274_ u2.mem\[53\]\[3\] _02486_ _02489_ u2.mem\[56\]\[3\] _02750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09013_ data_in_trans\[3\].data_sync _04134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06225_ _01577_ _01731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13005__CLK clknet_leaf_258_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08541__S _03836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06156_ _01617_ _01619_ _01663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11966__I _05971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10870__I _04986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06087_ _01556_ _01569_ _01593_ _01594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_104_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13155__CLK clknet_leaf_261_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09915_ _04707_ u2.mem\[41\]\[11\] _04701_ _04708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08340__I data_in_trans\[12\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09846_ _04573_ u2.mem\[40\]\[2\] _04661_ _04664_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08010__B1 _03459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09372__S _04358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09777_ _04624_ _00614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_06989_ _02410_ _02391_ _02424_ _02468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_39_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08728_ _03954_ _00235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_84_clock_I clknet_5_11_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08164__I1 u2.mem\[2\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08659_ _03909_ _00211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11206__I _05507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11670_ _04071_ _05769_ _05800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08716__S _03947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10621_ _05143_ _00939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13340_ _01219_ clknet_leaf_4_clock u2.mem\[160\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06627__B2 u2.mem\[161\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10552_ _05098_ _00915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13271_ _01150_ clknet_leaf_5_clock u2.mem\[148\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10483_ _05005_ u2.mem\[55\]\[5\] _05056_ _05058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09547__S _04474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12222_ _00101_ clknet_leaf_216_clock u2.mem\[6\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11223__I1 u2.mem\[151\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06035__I _01543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08451__S _03778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11876__I _05927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12153_ _00032_ clknet_leaf_56_clock u2.mem\[1\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10982__I0 _05343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11104_ _03487_ _05443_ _05444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_155_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12084_ output_active_hold\[2\] clknet_leaf_363_clock output_active_hold\[3\] vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_361_clock_I clknet_5_0_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12522__CLK clknet_leaf_112_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11035_ _05400_ _01096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06563__B1 _02047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11317__S _05576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10221__S _04887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12986_ _00865_ clknet_leaf_326_clock u2.mem\[53\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09352__I0 _04278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11937_ _05218_ u2.mem\[193\]\[10\] _05960_ _05963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06866__A1 _02339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08626__S _03885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11868_ _05922_ _01407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09104__I0 _04171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10819_ _05252_ _05263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__13028__CLK clknet_leaf_31_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11799_ _05880_ _01380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06618__A1 _02053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13538_ _01417_ clknet_leaf_34_clock u2.mem\[192\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06094__A2 _01600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07291__B2 u2.mem\[31\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13469_ _01348_ clknet_leaf_345_clock u2.mem\[181\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07830__A3 _03293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12052__CLK clknet_leaf_287_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06010_ u2.driver_mem\[1\] _01518_ _01519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__13178__CLK clknet_leaf_276_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07043__A1 _02429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07594__A2 _02906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07961_ _03421_ _03422_ _03423_ _03424_ _03425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_99_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09700_ _04565_ u2.mem\[37\]\[0\] _04567_ _04568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06912_ _02381_ _02391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_4_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07892_ u2.mem\[26\]\[13\] _02573_ _02575_ u2.mem\[10\]\[13\] _03358_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06149__A3 _01588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07346__A2 _02666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_106_clock_I clknet_5_11_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09631_ _04521_ _04527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_28_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06843_ _02319_ _02320_ _02321_ _02322_ _02323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_55_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11227__S _05520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_17_0_clock_I clknet_4_8_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09562_ _04157_ _04485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06774_ u2.mem\[168\]\[3\] _02093_ _02256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09343__I0 _04269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08513_ _03697_ _03820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09493_ _04440_ _04441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07649__A3 _03117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11150__I0 _05472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06857__A1 _02309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08444_ _03775_ _03776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_12_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08375_ _03734_ _00102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07326_ _02479_ _02801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08335__I data_in_trans\[11\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07282__A1 _02741_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06085__A2 _01591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07257_ u2.mem\[6\]\[2\] _02622_ _02624_ u2.mem\[47\]\[2\] _02734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06208_ _01714_ _01715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07188_ _02558_ _02666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12545__CLK clknet_leaf_168_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06139_ _01645_ _01646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06793__B1 _02088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08909__I0 _04044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10105__I _04819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10716__I0 _05198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12695__CLK clknet_leaf_110_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09582__I0 _04498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09829_ _04653_ _00637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12840_ _00719_ clknet_leaf_139_clock u2.mem\[44\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09334__I0 _04260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12771_ _00650_ clknet_leaf_90_clock u2.mem\[40\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11141__I0 _05466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11722_ _05831_ u2.mem\[182\]\[2\] _05827_ _05832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11653_ _05786_ u2.mem\[178\]\[0\] _05788_ _05789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_360_clock clknet_5_0_0_clock clknet_leaf_360_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_23_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12075__CLK clknet_2_2__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10604_ _05099_ u2.mem\[58\]\[2\] _05131_ _05134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11444__I1 u2.mem\[165\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11584_ _05719_ u2.mem\[173\]\[5\] _05738_ _05745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13320__CLK clknet_leaf_306_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13323_ _01202_ clknet_leaf_303_clock u2.mem\[157\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06076__A2 _01576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10535_ _05087_ _00909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13254_ _01133_ clknet_leaf_291_clock u2.mem\[145\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10466_ _05025_ u2.mem\[54\]\[14\] _05045_ _05048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12205_ _00084_ clknet_leaf_212_clock u2.mem\[5\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07025__A1 _02487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13185_ _01064_ clknet_leaf_277_clock u2.mem\[134\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13470__CLK clknet_leaf_347_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10397_ _04143_ _05004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07576__A2 _02890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12136_ _01462_ clknet_leaf_37_clock u2.driver_mem\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10015__I _04761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12067_ net22 clknet_2_1__leaf_clock_a data_in_trans\[9\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07328__A2 _02797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09573__I0 _04491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11018_ _05348_ _05390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11047__S _05404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06536__C2 u2.mem\[189\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_313_clock clknet_5_19_0_clock clknet_leaf_313_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09325__I0 _04246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07324__I _02476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12089__D net35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10886__S _05296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12969_ _00848_ clknet_leaf_125_clock u2.mem\[52\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06839__A1 u2.mem\[166\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06839__B2 u2.mem\[161\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06490_ u2.mem\[194\]\[14\] _01933_ _01977_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_328_clock clknet_5_7_0_clock clknet_leaf_328_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_92_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08160_ _03548_ u2.mem\[2\]\[1\] _03585_ _03587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08155__I _03582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07111_ _02577_ _02578_ _02463_ _02544_ _02590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__07264__A1 u2.mem\[27\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12568__CLK clknet_leaf_112_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08091_ _01980_ _03527_ _03536_ _00016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_32_clock_I clknet_5_3_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07042_ _02520_ _02521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10126__S _04835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10946__I0 _05343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07567__A2 _02881_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08993_ data_in_trans\[0\].data_sync _04117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07031__A4 _02468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06775__B1 _02086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06775__C2 _02088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07944_ _03405_ _03406_ _03407_ _03408_ _03409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_130_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09714__I _04138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_257_clock_I clknet_5_23_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06790__A3 _02250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07875_ _03337_ _03338_ _03339_ _03340_ _03341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_21_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11371__I0 _05591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09614_ _04517_ _00558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06826_ u2.mem\[164\]\[5\] _02051_ _02055_ u2.mem\[178\]\[5\] _02306_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09545_ _04139_ _04473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06757_ _01769_ _01996_ _02239_ _01476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12098__CLK clknet_leaf_224_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09476_ _04378_ u2.mem\[31\]\[9\] _04429_ _04431_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11674__I1 u2.mem\[179\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06688_ u2.mem\[151\]\[1\] _02085_ _02087_ u2.mem\[158\]\[1\] u2.mem\[193\]\[1\]
+ _02089_ _02172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_58_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13343__CLK clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08427_ _03698_ u2.mem\[7\]\[9\] _03764_ _03766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08358_ _03722_ _03723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08065__I data_in_trans\[8\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07309_ u2.mem\[32\]\[4\] _02782_ _02783_ u2.mem\[2\]\[4\] _02784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06058__A2 _01561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08289_ _03666_ _03667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09097__S _04192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10320_ _04955_ _00826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10251_ _04913_ u2.mem\[49\]\[12\] _04914_ _04915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10036__S _04777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10182_ _04864_ _04870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_132_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07191__B1 _02549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09560__S _04483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07730__A2 _03091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12823_ _00702_ clknet_leaf_135_clock u2.mem\[43\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11114__I0 _05430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_5_0_clock_I clknet_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08176__S _03595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12754_ _00633_ clknet_leaf_229_clock u2.mem\[39\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11665__I1 u2.mem\[178\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08530__I1 u2.mem\[9\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06916__C _02394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11705_ _05792_ u2.mem\[181\]\[2\] _05818_ _05821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12685_ _00564_ clknet_leaf_193_clock u2.mem\[35\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12710__CLK clknet_leaf_27_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11636_ _05285_ _05769_ _05778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11417__I1 u2.mem\[163\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08904__S _04061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07246__B2 u2.mem\[25\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11567_ _05735_ _01293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11330__S _05585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13306_ _01185_ clknet_leaf_358_clock u2.mem\[154\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10518_ _05072_ _05078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_116_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11498_ _05693_ _01266_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12860__CLK clknet_leaf_203_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13237_ _01116_ clknet_leaf_284_clock u2.mem\[143\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10449_ _05038_ _00872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09794__I0 _04605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06223__I _01572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13168_ _01047_ clknet_leaf_263_clock u2.mem\[131\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12119_ _01482_ clknet_leaf_332_clock u2.select_mem_col\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13099_ _00978_ clknet_leaf_245_clock u2.mem\[61\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10156__I1 u2.mem\[47\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_252_clock clknet_5_22_0_clock clknet_leaf_252_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11353__I0 _05589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07660_ _03122_ _03125_ _03128_ _03129_ _03130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_81_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07054__I _02532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12240__CLK clknet_leaf_227_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13366__CLK clknet_leaf_359_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07721__A2 _03072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06611_ _02064_ _02046_ _02096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07591_ _02555_ _03062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09330_ _04339_ _00452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11505__S _05691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06542_ _01988_ _02010_ _02027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11656__I1 u2.mem\[178\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_267_clock clknet_5_22_0_clock clknet_leaf_267_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_59_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09261_ _04298_ _00424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06473_ _01913_ _01964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12390__CLK clknet_leaf_77_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08212_ _03617_ _00056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09192_ _04251_ _04252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_159_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08143_ _03574_ _00030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11240__S _05529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08074_ _01962_ _03517_ _03524_ _00011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07025_ _02487_ _02496_ _02497_ _02434_ _02504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_134_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06460__A2 _01938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_205_clock clknet_5_29_0_clock clknet_leaf_205_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_162_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09645__S _04532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09785__I0 _04592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06133__I _01639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11592__I0 _05750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08976_ _04032_ u2.mem\[20\]\[8\] _04107_ _04108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input32_I mem_address_a[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09537__I0 _04467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07927_ u2.mem\[43\]\[14\] _03282_ _03283_ u2.mem\[20\]\[14\] _03392_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07858_ _02613_ _03325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07173__B1 _02489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07712__A2 _03170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06809_ _02286_ _02287_ _02288_ _02289_ _02290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_71_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07789_ u2.mem\[27\]\[12\] _03254_ _03255_ u2.mem\[35\]\[12\] _03256_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_77_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11415__S _05638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09528_ _04461_ _00528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_09459_ _04421_ _00499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06279__A2 _01782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07476__A1 u2.mem\[61\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11214__I _05513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12470_ _00349_ clknet_leaf_106_clock u2.mem\[21\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12883__CLK clknet_leaf_64_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11421_ _05633_ u2.mem\[163\]\[4\] _05637_ _05643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11150__S _05461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11352_ _05600_ _01213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08523__I _03799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10303_ _04889_ u2.mem\[51\]\[1\] _04944_ _04946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12113__CLK clknet_leaf_331_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_12_0_clock_I clknet_3_6_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11283_ _05557_ _01187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09776__I0 _04579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13022_ _00901_ clknet_leaf_259_clock u2.mem\[56\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10234_ _04902_ u2.mem\[49\]\[7\] _04896_ _04903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06043__I col_select_trans\[5\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06739__B1 _02089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10386__I1 u2.mem\[53\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06978__I _02456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10165_ _04815_ u2.mem\[47\]\[14\] _04856_ _04859_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12263__CLK clknet_leaf_55_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13389__CLK clknet_leaf_355_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07951__A2 _03246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10096_ _04819_ _04820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_47_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08200__I0 _03548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07164__B1 _02477_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09290__S _04313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07703__A2 _03114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11325__S _05575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12806_ _00685_ clknet_leaf_82_clock u2.mem\[42\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11638__I1 u2.mem\[177\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10998_ _05346_ u2.mem\[137\]\[3\] _05373_ _05377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07602__I _02586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09700__I0 _04565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07467__A1 u2.mem\[53\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12737_ _00616_ clknet_leaf_232_clock u2.mem\[38\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_205_clock_I clknet_5_29_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_9_0_clock_I clknet_3_4_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12668_ _00547_ clknet_leaf_193_clock u2.mem\[34\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07219__A1 u2.mem\[32\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08267__I0 _03572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07219__B2 u2.mem\[2\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11619_ _05767_ _01313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12599_ _00478_ clknet_leaf_113_clock u2.mem\[29\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11060__S _05413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10074__I0 _04804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08433__I _03753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06442__A2 _01924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07049__I _02527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09767__I0 _04565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12606__CLK clknet_leaf_195_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11574__I0 _05707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08830_ _03663_ _04017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09264__I _04289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_191_clock clknet_5_31_0_clock clknet_leaf_191_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_112_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08761_ _03962_ _03973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07712_ _03165_ _03170_ _03175_ _03180_ _03181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__12756__CLK clknet_leaf_69_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08692_ _03709_ _03932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08809__S _04000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07643_ u2.mem\[50\]\[9\] _03111_ _03112_ u2.mem\[51\]\[9\] _03113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07574_ _03037_ _03038_ _03041_ _03044_ _03045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_53_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09313_ _04278_ u2.mem\[27\]\[12\] _04328_ _04329_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07458__A1 u2.mem\[27\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06525_ row_select_trans\[3\].data_sync _02010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09244_ _04287_ _04288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_55_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06456_ _01945_ _01938_ _01947_ _01950_ _01470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06130__A1 u2.mem\[188\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06130__B2 u2.mem\[187\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12136__CLK clknet_leaf_37_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09175_ _04164_ u2.mem\[24\]\[11\] _04236_ _04240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08258__I0 _03563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10873__I _05296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06387_ u2.mem\[158\]\[5\] _01728_ _01729_ u2.mem\[151\]\[5\] _01577_ u2.mem\[193\]\[5\]
+ _01889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_147_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08126_ _03562_ _00025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08343__I _03659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_144_clock clknet_5_24_0_clock clknet_leaf_144_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_135_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06433__A2 _01931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08057_ _01878_ _03505_ _03512_ _00006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_162_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12286__CLK clknet_leaf_185_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07008_ _02346_ _02487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__06984__A3 _02382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10314__S _04949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_159_clock clknet_5_26_0_clock clknet_leaf_159_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_131_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06197__A1 _01552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07394__B1 _02867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08959_ _04098_ _00322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11317__I0 _05548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_1_clock_I clknet_5_0_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11209__I _03502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_154_clock_I clknet_5_27_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11970_ _05982_ _01449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07146__B1 _02624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10921_ _05326_ _05327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_3968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10852_ _05283_ _01030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07449__B2 u2.mem\[48\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10984__S _05365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13571_ _01450_ clknet_leaf_20_clock u2.mem\[194\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_10783_ _05213_ u2.mem\[62\]\[8\] _05242_ _05243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12522_ _00401_ clknet_leaf_112_clock u2.mem\[24\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06038__I _01544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06121__A1 u2.mem\[171\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06121__B2 u2.mem\[157\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08249__I0 _03554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12453_ _00332_ clknet_leaf_86_clock u2.mem\[20\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13061__CLK clknet_leaf_26_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06672__A2 _01999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_14_0_clock clknet_4_7_0_clock clknet_5_14_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_11404_ _05632_ _01233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12629__CLK clknet_leaf_97_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12384_ _00263_ clknet_leaf_221_clock u2.mem\[16\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07216__A4 _02693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_79_clock_I clknet_5_8_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11335_ _05507_ _05589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06424__A2 _01924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11266_ _05545_ _05546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_122_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10508__A1 _04224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10217_ _04572_ _04891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13005_ _00884_ clknet_leaf_258_clock u2.mem\[55\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12779__CLK clknet_leaf_253_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11197_ _04179_ _05482_ _05501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06188__A1 u2.mem\[146\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11181__A1 _04120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06188__B2 u2.mem\[186\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07924__A2 _02521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10148_ _04849_ _00760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10079_ _04601_ _04808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12009__CLK clknet_2_0__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09812__I _04638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06360__A1 u2.mem\[190\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06360__B2 u2.mem\[194\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07332__I _02488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08488__I0 _03802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10295__I0 _04918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06310_ _01810_ _01811_ _01812_ _01813_ _01814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__13404__CLK clknet_leaf_305_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_356_clock_I clknet_5_1_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07290_ u2.mem\[9\]\[3\] _02580_ _02582_ u2.mem\[25\]\[3\] _02766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06241_ u2.mem\[167\]\[1\] _01622_ _01623_ u2.mem\[183\]\[1\] _01747_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_61_clock clknet_5_9_0_clock clknet_leaf_61_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_106_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06172_ _01678_ _01644_ _01588_ _01679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_141_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13554__CLK clknet_leaf_14_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07000__C _02455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09931_ _04718_ _04719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_76_clock clknet_5_8_0_clock clknet_leaf_76_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_131_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11547__I0 _05711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09862_ _04596_ u2.mem\[40\]\[9\] _04671_ _04673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10134__S _04841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06179__A1 _01563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08813_ _03989_ _04005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_98_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09793_ _04617_ _04633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08744_ _03900_ u2.mem\[15\]\[0\] _03963_ _03964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08539__S _03836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09912__I0 _04705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08675_ _03920_ _00216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07679__B2 u2.mem\[24\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07626_ _03087_ _03090_ _03093_ _03096_ _03097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_96_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_14_clock clknet_5_3_0_clock clknet_leaf_14_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06351__A1 u2.mem\[145\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06351__B2 u2.mem\[163\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07557_ _02464_ _03028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13084__CLK clknet_leaf_261_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10286__I0 _04909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06508_ _01987_ _01991_ _01992_ _01993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_166_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07488_ u2.mem\[52\]\[6\] _02847_ _02848_ u2.mem\[21\]\[6\] _02961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06103__A1 _01607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07300__B1 _02614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09840__A2 _04659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_29_clock clknet_5_3_0_clock clknet_leaf_29_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09227_ _04163_ _04276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06439_ u2.mem\[193\]\[3\] _01928_ _01933_ u2.mem\[194\]\[3\] _01934_ _01937_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_155_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10038__I0 _04714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09158_ _04230_ _00389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_80_clock_I clknet_5_8_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08109_ _03550_ u2.mem\[1\]\[2\] _03546_ _03551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06406__A2 _01675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07603__B2 u2.mem\[31\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09089_ _04190_ _00360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12921__CLK clknet_leaf_159_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11120_ _05420_ u2.mem\[145\]\[0\] _05453_ _05454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11538__I0 _05717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11051_ _05392_ u2.mem\[140\]\[5\] _05403_ _05410_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07417__I _02527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10002_ _04716_ u2.mem\[43\]\[15\] _04755_ _04759_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07906__A2 _03369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09833__S _04654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08449__S _03778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06590__A1 _02007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11953_ _05903_ u2.mem\[194\]\[0\] _05972_ _05973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12301__CLK clknet_leaf_183_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13427__CLK clknet_leaf_349_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10904_ _05316_ _01049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08248__I _03634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06342__A1 u2.mem\[189\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11884_ _05933_ _01412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06342__B2 u2.mem\[180\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06893__A2 _02338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10835_ u2.mem\[63\]\[15\] _05229_ _05268_ _05272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10277__I0 _04900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13554_ _01433_ clknet_leaf_14_clock u2.mem\[193\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12451__CLK clknet_leaf_84_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10766_ _05233_ _00994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13577__CLK clknet_leaf_35_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12505_ _00384_ clknet_leaf_163_clock u2.mem\[23\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06645__A2 _02070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07842__B2 u2.mem\[22\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13485_ _01364_ clknet_leaf_289_clock u2.mem\[184\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10697_ _05117_ u2.mem\[60\]\[10\] _05184_ _05187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11402__I _05510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10029__I0 _04705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12436_ _00315_ clknet_leaf_107_clock u2.mem\[19\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_2_2__f_clock_a clknet_0_clock_a clknet_2_2__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08642__I0 _03829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12367_ _00246_ clknet_leaf_223_clock u2.mem\[15\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11318_ _05578_ _01201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12298_ _00177_ clknet_leaf_165_clock u2.mem\[10\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11529__I0 _05711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11249_ _05535_ _01175_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10201__I0 _04810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10889__S _05296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06790_ _02245_ _02249_ _02250_ _02271_ _02272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_110_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08359__S _03711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09542__I _04135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11701__I0 _05786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08460_ _03685_ u2.mem\[8\]\[6\] _03783_ _03786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06333__A1 u2.mem\[191\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07530__B1 _02914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06333__B2 u2.mem\[179\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07411_ u2.mem\[58\]\[5\] _02809_ _02810_ u2.mem\[36\]\[5\] _02885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08391_ _03727_ _03743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_23_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10268__I0 _04891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11513__S _05700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07342_ _02516_ _02817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07273_ u2.mem\[54\]\[3\] _02648_ _02649_ u2.mem\[55\]\[3\] _02749_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_102_clock_I clknet_5_11_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09012_ _04133_ _00340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12944__CLK clknet_leaf_235_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06224_ u2.mem\[163\]\[1\] _01643_ _01646_ u2.mem\[165\]\[1\] _01730_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11768__I0 _05831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06155_ u2.mem\[174\]\[0\] _01657_ _01659_ u2.mem\[155\]\[0\] _01661_ u2.mem\[181\]\[0\]
+ _01662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__08633__I0 _03820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07597__B1 _03067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08621__I _03879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06086_ _01573_ _01575_ _01593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_28_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09914_ _04601_ _04707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08010__A1 u2.active_mem\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09845_ _04663_ _00643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08010__B2 u2.active_mem\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12324__CLK clknet_leaf_84_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09776_ _04579_ u2.mem\[38\]\[4\] _04623_ _04624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_1543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_06988_ _02389_ _02467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_101_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_27_clock_I clknet_5_2_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08727_ _03926_ u2.mem\[14\]\[9\] _03952_ _03954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08658_ _03908_ u2.mem\[13\]\[1\] _03906_ _03909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12474__CLK clknet_leaf_123_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07609_ _02600_ _03080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08589_ _03815_ u2.mem\[11\]\[7\] _03862_ _03866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11423__S _05637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08077__A1 _01966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10620_ _05115_ u2.mem\[58\]\[9\] _05141_ _05143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10551_ _05097_ u2.mem\[57\]\[1\] _05095_ _05098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11222__I _05519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09828__S _04649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13270_ _01149_ clknet_leaf_5_clock u2.mem\[148\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10482_ _05057_ _00886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12221_ _00100_ clknet_leaf_213_clock u2.mem\[6\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08624__I0 _03811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12152_ _00031_ clknet_leaf_64_clock u2.mem\[1\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10431__I0 _05027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11103_ _05442_ _05443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_85_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_304_clock_I clknet_5_16_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12083_ output_active_hold\[1\] clknet_leaf_363_clock output_active_hold\[2\] vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09563__S _04483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11034_ _05390_ u2.mem\[139\]\[4\] _05394_ _05400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06051__I col_select_trans\[2\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06986__I _02464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06563__A1 u2.mem\[180\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09362__I _04357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06563__B2 u2.mem\[150\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12985_ _00864_ clknet_leaf_319_clock u2.mem\[53\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11936_ _05962_ _01435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08907__S _04066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06866__A2 _02344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11867_ _05911_ u2.mem\[191\]\[3\] _05918_ _05922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06935__B _02411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09104__I1 u2.mem\[22\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12967__CLK clknet_leaf_124_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11333__S _05585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08068__A1 _01954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08706__I _03941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10818_ _05262_ _01017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07610__I _02602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11798_ _05864_ u2.mem\[187\]\[0\] _05879_ _05880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06618__A2 _02012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13537_ _01416_ clknet_leaf_14_clock u2.mem\[192\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08863__I0 _04039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10749_ _05221_ _00989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11132__I _05334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09738__S _04593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10670__I0 _05128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06226__I _01589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07291__A2 _02585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13468_ _01347_ clknet_leaf_346_clock u2.mem\[181\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11991__CLK clknet_leaf_318_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12419_ _00298_ clknet_leaf_110_clock u2.mem\[18\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08615__I0 _03802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13399_ _01278_ clknet_leaf_297_clock u2.mem\[170\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10422__I0 _05020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07043__A2 _02445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12347__CLK clknet_leaf_221_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06251__B1 _01631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07960_ u2.mem\[3\]\[15\] _03267_ _02358_ _03424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06911_ _02389_ _02390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__09040__I0 _04154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07891_ _03353_ _03354_ _03355_ _03356_ _03357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_68_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09630_ _04526_ _00565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10412__S _05012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06842_ u2.mem\[145\]\[5\] _02082_ _02094_ u2.mem\[168\]\[5\] _02322_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12497__CLK clknet_leaf_163_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07751__B1 _03121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09561_ _04484_ _00538_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06773_ _02251_ _02252_ _02253_ _02254_ _02255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_167_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08512_ _03819_ _00154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10211__I _04886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06306__A1 u2.mem\[178\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09492_ _03478_ _03986_ _04439_ _04440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_93_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06306__B2 u2.mem\[164\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11150__I1 u2.mem\[146\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06857__A2 _02314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08443_ mem_address_trans\[2\].data_sync _03774_ _03775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08374_ _03676_ u2.mem\[6\]\[4\] _03733_ _03734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08059__A1 _03513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07325_ u2.mem\[16\]\[4\] _02798_ _02799_ u2.mem\[33\]\[4\] _02800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08854__I0 _04032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_253_clock_I clknet_5_22_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07256_ u2.mem\[8\]\[2\] _02612_ _02614_ u2.mem\[4\]\[2\] _02733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10661__I0 _05119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06136__I _01642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06085__A3 _01588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13122__CLK clknet_leaf_242_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06207_ _01557_ _01619_ _01714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07187_ _02639_ _02644_ _02653_ _02664_ _02665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_105_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06138_ _01570_ _01644_ _01600_ _01645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_30_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08351__I data_in_trans\[14\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07034__A2 _02501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06242__B1 _01614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13272__CLK clknet_5_0_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06069_ _01573_ _01575_ _01549_ _01576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__11118__A1 _05285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06793__B2 u2.mem\[193\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09031__I0 _04148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09828_ _04602_ u2.mem\[39\]\[11\] _04649_ _04653_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07742__B1 _03032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09759_ _04612_ u2.mem\[37\]\[14\] _04606_ _04613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11217__I _03510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09334__I1 u2.mem\[28\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12770_ _00649_ clknet_leaf_155_clock u2.mem\[40\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11141__I1 u2.mem\[146\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11721_ _03666_ _05831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08526__I _03714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11652_ _05787_ _05788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_39_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06474__C _01964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10603_ _05133_ _00931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10992__S _05373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11583_ _05744_ _01300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13322_ _01201_ clknet_leaf_342_clock u2.mem\[157\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10652__I0 _05110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08462__S _03783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10534_ _05018_ u2.mem\[56\]\[11\] _05083_ _05087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07273__A2 _02648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10791__I _05231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13253_ _01132_ clknet_leaf_291_clock u2.mem\[145\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10465_ _05047_ _00879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12204_ _00083_ clknet_leaf_211_clock u2.mem\[5\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13184_ _01063_ clknet_leaf_277_clock u2.mem\[134\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10396_ _05003_ _00854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12135_ _01461_ clknet_leaf_37_clock u2.driver_mem\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06784__A1 u2.mem\[170\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06784__B2 u2.mem\[156\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09022__I0 _04140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12066_ data_in_trans\[8\].A clknet_leaf_32_clock data_in_trans\[8\].data_sync vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11017_ _05389_ _01089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06536__A1 u2.mem\[176\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09092__I _04181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06536__B2 u2.mem\[172\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12968_ _00847_ clknet_leaf_124_clock u2.mem\[52\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08637__S _03890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11919_ _05909_ u2.mem\[193\]\[2\] _05950_ _05953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12899_ _00778_ clknet_leaf_64_clock u2.mem\[48\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13145__CLK clknet_leaf_39_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07110_ _02571_ _02576_ _02583_ _02588_ _02589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_147_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10643__I0 _05101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08090_ _03535_ _03529_ _03536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07264__A2 _02428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11797__I _05878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07041_ _02394_ _02438_ _02439_ _02519_ _02520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_31_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11199__I1 u2.mem\[150\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06224__B1 _01646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08992_ _04116_ _00337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06775__A1 u2.mem\[151\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06775__B2 u2.mem\[158\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07943_ u2.mem\[18\]\[14\] _03316_ _03317_ u2.mem\[19\]\[14\] _03408_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_1313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11238__S _05529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07874_ u2.mem\[3\]\[13\] _03267_ _03211_ _03340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07724__B1 _03078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11371__I1 u2.mem\[160\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09613_ _04491_ u2.mem\[34\]\[12\] _04516_ _04517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06825_ u2.mem\[171\]\[5\] _02066_ _02068_ u2.mem\[157\]\[5\] _02305_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09544_ _04472_ _00533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06756_ _02209_ _02214_ _02223_ _02238_ _02239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_83_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10876__I _04991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09475_ _04430_ _00506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06687_ _02164_ _02165_ _02166_ _02170_ _02171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_34_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08426_ _03765_ _00122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08346__I data_in_trans\[13\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08357_ _03721_ _03722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12512__CLK clknet_leaf_162_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11587__A1 _04393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07308_ _02395_ _02783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07255__A2 _02617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08288_ _03499_ _03666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07239_ u2.mem\[61\]\[2\] _02666_ _02667_ u2.mem\[63\]\[2\] _02716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09177__I _04225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10250_ _04886_ _04914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_133_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10181_ _04869_ _00773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09905__I _04682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07963__B1 _02511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13018__CLK clknet_leaf_322_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06518__A1 _02000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07425__I _02558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12822_ _00701_ clknet_leaf_83_clock u2.mem\[43\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12042__CLK clknet_leaf_299_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13168__CLK clknet_leaf_263_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09640__I _04521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11114__I1 u2.mem\[144\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12753_ _00632_ clknet_leaf_230_clock u2.mem\[39\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11704_ _05820_ _01345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12684_ _00563_ clknet_leaf_193_clock u2.mem\[35\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08818__I0 _03937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12192__CLK clknet_leaf_228_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11635_ _05777_ _01319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09288__S _04313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07246__A2 _02580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11566_ _05715_ u2.mem\[172\]\[3\] _05731_ _05735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_149_clock_I clknet_5_24_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13305_ _01184_ clknet_leaf_358_clock u2.mem\[154\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10517_ _05077_ _00901_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11497_ _05663_ u2.mem\[168\]\[0\] _05692_ _05693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13236_ _01115_ clknet_leaf_273_clock u2.mem\[142\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06504__I row_select_trans\[3\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10448_ _05007_ u2.mem\[54\]\[6\] _05035_ _05038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13167_ _01046_ clknet_leaf_263_clock u2.mem\[131\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06757__A1 _01769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10379_ _04990_ _00850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12118_ _01481_ clknet_leaf_334_clock u2.select_mem_col\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_201_clock_I clknet_5_28_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13098_ _00977_ clknet_leaf_45_clock u2.mem\[60\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11058__S _05413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12049_ net7 clknet_2_3__leaf_clock_a data_in_trans\[0\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07335__I _02499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11353__I1 u2.mem\[159\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10897__S _05310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06610_ u2.mem\[177\]\[0\] _02092_ _02094_ u2.mem\[168\]\[0\] _02095_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_94_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07590_ _02553_ _03061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08367__S _03728_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06541_ _02016_ _02025_ _02026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12535__CLK clknet_leaf_115_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09260_ _04265_ u2.mem\[26\]\[6\] _04295_ _04298_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08166__I _03584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10864__I0 _05202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06472_ u2.mem\[194\]\[10\] _01946_ _01963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07070__I _02548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08211_ _03559_ u2.mem\[3\]\[6\] _03614_ _03617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09191_ _04249_ _04250_ _04251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08809__I0 _03928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08142_ _03572_ u2.mem\[1\]\[12\] _03573_ _03574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12685__CLK clknet_leaf_193_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08073_ _03523_ _03519_ _03524_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07024_ _02502_ _02503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06414__I _01914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11041__I0 _05380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06748__A1 u2.mem\[154\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07945__B1 _02629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11592__I1 u2.mem\[174\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06748__B2 u2.mem\[162\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06212__A3 _01596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08975_ _04096_ _04107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_9_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07926_ u2.mem\[49\]\[14\] _02531_ _02533_ u2.mem\[46\]\[14\] _03391_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12065__CLK clknet_2_3__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09661__S _04544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input25_I mem_address_a[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13310__CLK clknet_leaf_348_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07857_ _02611_ _03324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07173__A1 u2.mem\[53\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07173__B2 u2.mem\[56\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07712__A3 _03175_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06808_ u2.mem\[155\]\[4\] _02030_ _02192_ u2.mem\[150\]\[4\] _02289_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10600__S _05131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07788_ _02435_ _03255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09527_ _04389_ u2.mem\[32\]\[14\] _04458_ _04461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06739_ u2.mem\[177\]\[2\] _02092_ _02089_ u2.mem\[193\]\[2\] _02222_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_09458_ _04360_ u2.mem\[31\]\[1\] _04419_ _04421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07476__A2 _02899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08409_ _03664_ u2.mem\[7\]\[1\] _03754_ _03756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09389_ _04375_ u2.mem\[29\]\[8\] _04376_ _04377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11420_ _05642_ _01239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08804__I _03989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07228__A2 _02645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_150_clock_I clknet_5_25_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06436__B1 _01933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11351_ _05587_ u2.mem\[159\]\[1\] _05598_ _05600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_312_clock clknet_5_17_0_clock clknet_leaf_312_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10302_ _04945_ _00818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09225__I0 _04274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11282_ _05556_ u2.mem\[154\]\[5\] _05545_ _05557_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11032__I0 _05388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13021_ _00900_ clknet_leaf_258_clock u2.mem\[56\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10233_ _04588_ _04902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06739__A1 u2.mem\[177\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06739__B2 u2.mem\[193\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10164_ _04858_ _00767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_327_clock clknet_5_7_0_clock clknet_leaf_327_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_43_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10095_ _04394_ _04760_ _04819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_120_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07155__I _02443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10299__A1 _04072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_10_0_clock clknet_4_5_0_clock clknet_5_10_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_78_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_75_clock_I clknet_5_8_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06994__I _02412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10510__S _05073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08187__S _03600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12805_ _00684_ clknet_leaf_82_clock u2.mem\[42\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10997_ _05376_ _01082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11405__I _05513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12736_ _00615_ clknet_leaf_229_clock u2.mem\[38\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09700__I1 u2.mem\[37\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12667_ _00546_ clknet_leaf_195_clock u2.mem\[34\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11618_ _05758_ u2.mem\[175\]\[5\] _05760_ _05767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08267__I1 u2.mem\[4\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12598_ _00477_ clknet_leaf_96_clock u2.mem\[29\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11549_ _05713_ u2.mem\[171\]\[2\] _05722_ _05725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11140__I _05342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09746__S _04593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09767__I1 u2.mem\[38\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13219_ _01098_ clknet_leaf_283_clock u2.mem\[140\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12088__CLK clknet_leaf_298_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09545__I _04139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11574__I1 u2.mem\[173\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13333__CLK clknet_leaf_4_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_352_clock_I clknet_5_1_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08760_ _03972_ _00249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07065__I _02347_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07711_ _03176_ _03177_ _03178_ _03179_ _03180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08691_ _03931_ _00221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13483__CLK clknet_leaf_290_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07642_ _02504_ _03112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07573_ u2.mem\[58\]\[8\] _03042_ _03043_ u2.mem\[36\]\[8\] _03044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09312_ _04312_ _04328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_40_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06524_ _02008_ _02009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09243_ _03581_ _04247_ _04287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_166_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06455_ u2.mem\[193\]\[6\] _01942_ _01948_ u2.mem\[192\]\[6\] _01949_ _01950_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06130__A2 _01631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09174_ _04239_ _00396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08258__I1 u2.mem\[4\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06386_ u2.mem\[177\]\[5\] _01583_ _01646_ u2.mem\[165\]\[5\] u2.mem\[163\]\[5\]
+ _01642_ _01888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_108_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08125_ _03561_ u2.mem\[1\]\[7\] _03555_ _03562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11262__I0 _05517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08056_ _03511_ _03508_ _03512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07007_ _02485_ _02486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11714__A1 _04179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09455__I _04418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06197__A2 _01615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07394__B2 u2.mem\[34\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08958_ _04010_ u2.mem\[20\]\[0\] _04097_ _04098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12700__CLK clknet_leaf_256_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11317__I1 u2.mem\[157\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07909_ u2.mem\[45\]\[14\] _02444_ _02448_ u2.mem\[34\]\[14\] _03374_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_3914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08889_ _04023_ u2.mem\[18\]\[4\] _04056_ _04057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10330__S _04959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10920_ _04121_ _05317_ _05326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_72_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09190__I _03987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12850__CLK clknet_leaf_150_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10851_ _05204_ u2.mem\[128\]\[4\] _05277_ _05283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13570_ _01449_ clknet_leaf_14_clock u2.mem\[194\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09694__I0 _04498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10782_ _05231_ _05242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_12521_ _00400_ clknet_leaf_118_clock u2.mem\[24\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13206__CLK clknet_leaf_271_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_12452_ _00331_ clknet_leaf_84_clock u2.mem\[20\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09446__I0 _04387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_251_clock clknet_5_22_0_clock clknet_leaf_251_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11403_ _05631_ u2.mem\[162\]\[3\] _05625_ _05632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12383_ _00262_ clknet_leaf_223_clock u2.mem\[16\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09566__S _04483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12230__CLK clknet_leaf_69_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11334_ _05588_ _01207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13356__CLK clknet_leaf_360_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11265_ _04287_ _05527_ _05545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__10505__S _05066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09365__I _04127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07909__B1 _02448_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_266_clock clknet_5_23_0_clock clknet_leaf_266_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13004_ _00883_ clknet_leaf_257_clock u2.mem\[55\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10216_ _04890_ _00787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11196_ _05499_ _05500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07385__A1 u2.mem\[8\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12380__CLK clknet_leaf_205_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11181__A2 _05482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10147_ _04797_ u2.mem\[47\]\[6\] _04846_ _04849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10078_ _04807_ _00732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07137__A1 _02568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08185__I0 _03572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11336__S _05585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07688__A2 _03094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07613__I _02607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_204_clock clknet_5_29_0_clock clknet_leaf_204_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_22_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_1551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09685__I0 _04489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08101__A3 _03544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11492__I0 _05680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12719_ _00598_ clknet_leaf_236_clock u2.mem\[37\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11071__S _05422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06240_ u2.mem\[178\]\[1\] _01618_ _01620_ u2.mem\[164\]\[1\] _01746_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09437__I0 _04378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_219_clock clknet_5_28_0_clock clknet_leaf_219_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_102_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06171_ _01677_ _01678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_129_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08380__S _03733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09930_ _04288_ _04659_ _04718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06899__I _02377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10415__S _05012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12723__CLK clknet_leaf_71_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11547__I1 u2.mem\[171\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09861_ _04672_ _00650_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06179__A2 _01677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08812_ _04004_ _00269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09792_ _04632_ _00621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08743_ _03962_ _03963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08176__I0 _03563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07128__A1 _02466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11246__S _05528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07679__A2 _03077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08674_ _03919_ u2.mem\[13\]\[6\] _03915_ _03920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07625_ u2.mem\[6\]\[8\] _03094_ _03095_ u2.mem\[47\]\[8\] _03096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13229__CLK clknet_leaf_286_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06351__A2 _01639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07556_ u2.mem\[15\]\[8\] _03025_ _03026_ u2.mem\[13\]\[8\] _03027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06139__I _01645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08555__S _03846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09676__I0 _04480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06507_ row_select_trans\[5\].data_sync row_select_trans\[4\].data_sync _01992_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07487_ u2.mem\[17\]\[6\] _02844_ _02845_ u2.mem\[24\]\[6\] _02960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06103__A2 _01609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09226_ _04275_ _00412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09428__I0 _04369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12253__CLK clknet_leaf_213_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06438_ u2.mem\[192\]\[3\] _01931_ _01936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09157_ _04136_ u2.mem\[24\]\[3\] _04226_ _04230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06369_ u2.mem\[146\]\[4\] _01691_ _01693_ u2.mem\[186\]\[4\] _01872_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_23_clock_I clknet_5_2_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08108_ _03500_ _03550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07064__B1 _02542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07603__A2 _03072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09088_ _04148_ u2.mem\[22\]\[6\] _04187_ _04190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08039_ _01727_ _03490_ _03498_ _00002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_150_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10325__S _04954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11050_ _05409_ _01102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06602__I _02086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10001_ _04758_ _00704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07906__A3 _03370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_248_clock_I clknet_5_22_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08167__I0 _03554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06590__A2 _02037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08529__I _03718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11952_ _05971_ _05972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_123_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07433__I _02574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10903_ _05307_ u2.mem\[131\]\[5\] _05309_ _05316_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11883_ u2.mem\[192\]\[2\] _03500_ _05932_ _05933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10834_ _05271_ _01024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08465__S _03788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09667__I0 _04471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06893__A3 _02344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_300_clock_I clknet_5_17_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11474__I0 _05677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13553_ _01432_ clknet_leaf_14_clock u2.mem\[193\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10765_ _05194_ u2.mem\[62\]\[0\] _05232_ _05233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12504_ _00383_ clknet_leaf_121_clock u2.mem\[23\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_190_clock clknet_5_31_0_clock clknet_leaf_190_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_73_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07842__A2 _03146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09419__I0 _04360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13484_ _01363_ clknet_leaf_290_clock u2.mem\[184\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10696_ _05186_ _00971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10029__I1 u2.mem\[44\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12435_ _00314_ clknet_leaf_108_clock u2.mem\[19\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12746__CLK clknet_leaf_50_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07055__B1 _02533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12366_ _00245_ clknet_leaf_209_clock u2.mem\[15\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08642__I1 u2.mem\[12\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11317_ _05548_ u2.mem\[157\]\[1\] _05576_ _05578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06802__C2 u2.mem\[192\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12297_ _00176_ clknet_leaf_120_clock u2.mem\[10\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11529__I1 u2.mem\[170\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06512__I row_select_trans\[4\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12896__CLK clknet_leaf_224_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11248_ _05517_ u2.mem\[152\]\[5\] _05528_ _05535_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11179_ _05472_ u2.mem\[148\]\[5\] _05483_ _05490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08158__I0 _03539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11066__S _05412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11701__I1 u2.mem\[181\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_143_clock clknet_5_24_0_clock clknet_leaf_143_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_97_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07530__B2 u2.mem\[22\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07410_ u2.mem\[53\]\[5\] _02806_ _02807_ u2.mem\[56\]\[5\] _02884_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12276__CLK clknet_leaf_102_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08390_ _03742_ _00109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13521__CLK clknet_leaf_16_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07341_ _02514_ _02816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_158_clock clknet_5_26_0_clock clknet_leaf_158_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_32_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07294__B1 _02593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07272_ u2.mem\[50\]\[3\] _02645_ _02646_ u2.mem\[51\]\[3\] _02748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09011_ _04132_ u2.mem\[21\]\[2\] _04124_ _04133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06223_ _01572_ _01729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11768__I1 u2.mem\[185\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06154_ _01660_ _01661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_197_clock_I clknet_5_30_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08633__I1 u2.mem\[12\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06085_ _01564_ _01591_ _01588_ _01592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__09934__S _04719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09913_ _04706_ _00668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09844_ _04570_ u2.mem\[40\]\[1\] _04661_ _04663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08010__A2 _03458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09733__I _04566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06021__A1 u2.driver_mem\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09775_ _04617_ _04623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_41_1533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10879__I _04994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_06987_ _02387_ _02466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_3018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13051__CLK clknet_leaf_254_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08726_ _03953_ _00234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08657_ _03663_ _03908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07608_ u2.mem\[17\]\[8\] _03077_ _03078_ u2.mem\[24\]\[8\] _03079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08588_ _03865_ _00184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07539_ _03007_ _03008_ _03009_ _03010_ _03011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_23_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08077__A2 _03517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12769__CLK clknet_leaf_154_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10550_ _04991_ _05097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07285__B1 _02542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09209_ _04263_ u2.mem\[25\]\[5\] _04261_ _04264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10481_ _05001_ u2.mem\[55\]\[4\] _05056_ _05057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12220_ _00099_ clknet_leaf_215_clock u2.mem\[6\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08624__I1 u2.mem\[12\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12151_ _00030_ clknet_leaf_64_clock u2.mem\[1\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10431__I1 u2.mem\[53\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09844__S _04661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11102_ _03984_ _03985_ _05274_ _05442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_150_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12082_ output_active_hold\[0\] clknet_leaf_363_clock output_active_hold\[1\] vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12149__CLK clknet_leaf_73_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11033_ _05399_ _01095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_60_clock clknet_5_12_0_clock clknet_leaf_60_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_18_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12299__CLK clknet_leaf_170_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12984_ _00863_ clknet_leaf_329_clock u2.mem\[53\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13544__CLK clknet_leaf_32_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11695__I0 _05796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11935_ _05216_ u2.mem\[193\]\[9\] _05960_ _05962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07512__A1 u2.mem\[58\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11614__S _05761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11866_ _05921_ _01406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_75_clock clknet_5_8_0_clock clknet_leaf_75_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_33_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06935__C _02413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10817_ u2.mem\[63\]\[7\] _03515_ _05258_ _05262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08068__A2 _03517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11797_ _05878_ _05879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08312__I0 _03685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13536_ _01415_ clknet_leaf_318_clock u2.mem\[192\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08923__S _04074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10748_ _05220_ u2.mem\[61\]\[11\] _05214_ _05221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13467_ _01346_ clknet_leaf_346_clock u2.mem\[181\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10679_ _05099_ u2.mem\[60\]\[2\] _05174_ _05177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12418_ _00297_ clknet_leaf_160_clock u2.mem\[18\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13398_ _01277_ clknet_leaf_307_clock u2.mem\[169\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12349_ _00228_ clknet_leaf_202_clock u2.mem\[14\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07043__A3 _02446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_13_clock clknet_5_3_0_clock clknet_leaf_13_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_86_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06251__B2 u2.mem\[188\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13074__CLK clknet_leaf_241_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06910_ _02366_ _02367_ _02368_ _02389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_4_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07890_ u2.mem\[57\]\[13\] _03294_ _03295_ u2.mem\[41\]\[13\] _03356_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07200__B1 _02587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06841_ u2.mem\[151\]\[5\] _02085_ _02087_ u2.mem\[158\]\[5\] u2.mem\[193\]\[5\]
+ _02089_ _02321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_67_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_28_clock clknet_5_3_0_clock clknet_leaf_28_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_3_1313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09560_ _04482_ u2.mem\[33\]\[8\] _04483_ _04484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06772_ u2.mem\[184\]\[3\] _02072_ _01994_ _02254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08511_ _03817_ u2.mem\[9\]\[8\] _03818_ _03819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09491_ _03984_ _03985_ _04439_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12911__CLK clknet_leaf_157_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08442_ mem_address_trans\[3\].data_sync _03774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_169_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06857__A3 _02323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06711__C1 _02127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11438__I0 _05635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08373_ _03727_ _03733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_56_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07324_ _02476_ _02799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07267__B1 _02471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10110__I0 _04797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07255_ u2.mem\[39\]\[2\] _02617_ _02619_ u2.mem\[48\]\[2\] _02732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07282__A3 _02752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09728__I _04588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06206_ _01712_ _01713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07186_ _02656_ _02659_ _02662_ _02663_ _02664_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_145_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11610__I0 _05750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06137_ _01593_ _01644_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13417__CLK clknet_leaf_298_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06242__A1 u2.mem\[171\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06152__I _01658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06242__B2 u2.mem\[157\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06068_ _01574_ _01575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__11118__A2 _05443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06793__A2 _02091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07990__B2 u2.mem\[4\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09031__I1 u2.mem\[21\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12441__CLK clknet_leaf_127_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09827_ _04652_ _00636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13567__CLK clknet_leaf_15_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09758_ _04611_ _04612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08079__I data_in_trans\[12\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08709_ _03908_ u2.mem\[14\]\[1\] _03942_ _03944_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09689_ _04560_ _00590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12591__CLK clknet_leaf_172_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11720_ _05830_ _01351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11651_ _05295_ _05769_ _05787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_14_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11054__A1 _05411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10602_ _05097_ u2.mem\[58\]\[1\] _05131_ _05133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10101__I0 _04788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11582_ _05717_ u2.mem\[173\]\[4\] _05738_ _05744_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13321_ _01200_ clknet_leaf_303_clock u2.mem\[157\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10533_ _05086_ _00908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13252_ _01131_ clknet_leaf_291_clock u2.mem\[145\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10464_ _05023_ u2.mem\[54\]\[13\] _05045_ _05047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12203_ _00082_ clknet_leaf_217_clock u2.mem\[5\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11601__I0 _05756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13183_ _01062_ clknet_leaf_273_clock u2.mem\[134\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10395_ _05001_ u2.mem\[53\]\[4\] _05002_ _05003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06233__A1 u2.mem\[173\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06233__B2 u2.mem\[185\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12134_ _01460_ clknet_leaf_14_clock u2.driver_mem\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12065_ net21 clknet_2_3__leaf_clock_a data_in_trans\[8\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09022__I1 u2.mem\[21\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11016_ _05388_ u2.mem\[138\]\[3\] _05382_ _05389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07733__A1 _03186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11408__I _05516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07107__B _02453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12934__CLK clknet_leaf_31_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_145_clock_I clknet_5_24_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11668__I0 _05798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12967_ _00846_ clknet_leaf_124_clock u2.mem\[52\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08533__I0 _03833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07497__B1 _02948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11918_ _05952_ _01427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12898_ _00777_ clknet_leaf_230_clock u2.mem\[48\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07621__I _02613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11849_ _05910_ _01400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11143__I _05345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07249__B1 _02681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12314__CLK clknet_leaf_118_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13519_ _01398_ clknet_leaf_16_clock u2.mem\[190\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07040_ _02410_ _02403_ _02383_ _02519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_62_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07068__I _02347_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06224__A1 u2.mem\[163\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12464__CLK clknet_leaf_173_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07421__B1 _02894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06224__B2 u2.mem\[165\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08991_ _04048_ u2.mem\[20\]\[15\] _04112_ _04116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07972__A1 _03420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06775__A2 _02084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07942_ u2.mem\[52\]\[14\] _03313_ _03314_ u2.mem\[21\]\[14\] _03407_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09283__I _04310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07873_ u2.mem\[16\]\[13\] _03264_ _03265_ u2.mem\[33\]\[13\] _03339_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09612_ _04500_ _04516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_83_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06824_ _01844_ _01996_ _02304_ _01478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08828__S _04015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09543_ _04471_ u2.mem\[33\]\[3\] _04465_ _04472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11659__I0 _05792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06755_ _02224_ _02231_ _02232_ _02237_ _02238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_43_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08524__I0 _03826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11254__S _05537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11284__A1 _04310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09474_ _04375_ u2.mem\[31\]\[8\] _04429_ _04430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06686_ u2.mem\[146\]\[1\] _02156_ _02158_ u2.mem\[186\]\[1\] _02169_ _02170_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08425_ _03693_ u2.mem\[7\]\[8\] _03764_ _03765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_347_clock_I clknet_5_4_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06147__I _01653_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08356_ data_in_trans\[15\].data_sync _03721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07307_ _02385_ _02782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11587__A2 _05729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11831__I0 _05870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10892__I _05309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08287_ _03665_ _00083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07238_ _02699_ _02704_ _02709_ _02714_ _02715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_30_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12807__CLK clknet_leaf_140_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07169_ u2.mem\[50\]\[1\] _02645_ _02646_ u2.mem\[51\]\[1\] _02647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10180_ _04790_ u2.mem\[48\]\[3\] _04865_ _04869_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12957__CLK clknet_leaf_196_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06518__A2 _02002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10570__I0 _05110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07191__A2 _02546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12821_ _00700_ clknet_leaf_83_clock u2.mem\[43\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11164__S _05474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12752_ _00631_ clknet_leaf_227_clock u2.mem\[39\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11703_ _05790_ u2.mem\[181\]\[1\] _05818_ _05820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12683_ _00562_ clknet_leaf_195_clock u2.mem\[35\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12337__CLK clknet_leaf_152_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09569__S _04483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11634_ _05758_ u2.mem\[176\]\[5\] _05770_ _05777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06057__I _01563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11565_ _05734_ _01292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09368__I _04131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13304_ _01183_ clknet_leaf_362_clock u2.mem\[154\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12487__CLK clknet_leaf_121_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10516_ _04998_ u2.mem\[56\]\[3\] _05073_ _05077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11496_ _05691_ _05692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_143_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_71_clock_I clknet_5_8_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13235_ _01114_ clknet_leaf_272_clock u2.mem\[142\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10447_ _05037_ _00871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13166_ _01045_ clknet_leaf_263_clock u2.mem\[131\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10378_ _04987_ u2.mem\[53\]\[0\] _04989_ _04990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11339__S _05585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07954__B2 u2.mem\[30\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12117_ _01480_ clknet_leaf_332_clock u2.select_mem_col\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13097_ _00976_ clknet_leaf_45_clock u2.mem\[60\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12048_ col_select_trans\[5\].A clknet_leaf_288_clock col_select_trans\[5\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__06520__I row_select_trans\[5\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11889__I0 u2.mem\[192\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_296_clock_I clknet_5_17_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10561__I0 _05103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13112__CLK clknet_leaf_39_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10977__I _05364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06390__B1 _01630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11074__S _05422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06540_ _02024_ _02025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07351__I _02541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06471_ u2.mem\[0\]\[10\] _01962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13262__CLK clknet_leaf_271_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08210_ _03616_ _00055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11802__S _05879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09190_ _03987_ _04250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08383__S _03738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08141_ _03545_ _03573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_119_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11813__I0 _05864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10418__S _05012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06445__A1 u2.mem\[192\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08072_ data_in_trans\[10\].data_sync _03523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07023_ _02483_ _02491_ _02492_ _02393_ _02502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_134_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08974_ _04106_ _00329_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07925_ u2.mem\[14\]\[14\] _02526_ _02528_ u2.mem\[12\]\[14\] _03390_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_151_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09698__A1 _04121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07856_ u2.mem\[39\]\[12\] _03321_ _03322_ u2.mem\[48\]\[12\] _03323_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07173__A2 _02486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06807_ u2.mem\[174\]\[4\] _02035_ _02039_ u2.mem\[181\]\[4\] _02288_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input18_I data_in_a[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07787_ _02427_ _03254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09526_ _04460_ _00527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06738_ u2.mem\[151\]\[2\] _02085_ _02087_ u2.mem\[158\]\[2\] u2.mem\[168\]\[2\]
+ _02094_ _02221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_101_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09457_ _04420_ _00498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06669_ u2.mem\[179\]\[0\] _02151_ _02153_ u2.mem\[191\]\[0\] _02154_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09389__S _04376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08408_ _03755_ _00114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06684__A1 u2.mem\[179\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09388_ _04357_ _04376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07881__B1 _02523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06684__B2 u2.mem\[191\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08339_ _03707_ _00093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11804__I0 _05872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10328__S _04959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06436__A1 u2.mem\[193\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11350_ _05599_ _01212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06436__B2 u2.mem\[194\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10301_ _04885_ u2.mem\[51\]\[0\] _04944_ _04945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11281_ _05516_ _05556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09225__I1 u2.mem\[25\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13020_ _00899_ clknet_leaf_258_clock u2.mem\[56\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10232_ _04901_ _00792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06739__A2 _02092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10163_ _04813_ u2.mem\[47\]\[13\] _04856_ _04858_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13135__CLK clknet_leaf_314_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10094_ _04818_ _00737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10998__S _05373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08736__I0 _03935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10299__A2 _04863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10543__I0 _05027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07164__A2 _02475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_18_clock_I clknet_5_2_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13285__CLK clknet_leaf_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12804_ _00683_ clknet_leaf_62_clock u2.mem\[42\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10996_ _05343_ u2.mem\[137\]\[2\] _05373_ _05376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07171__I _02510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12735_ _00614_ clknet_leaf_237_clock u2.mem\[38\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12666_ _00545_ clknet_leaf_56_clock u2.mem\[33\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11617_ _05766_ _01312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10238__S _04905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12597_ _00476_ clknet_leaf_99_clock u2.mem\[29\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11548_ _05724_ _01285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06515__I _01999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11479_ _05681_ _01259_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13218_ _01097_ clknet_leaf_283_clock u2.mem\[139\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07927__B2 u2.mem\[20\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13149_ _01028_ clknet_leaf_264_clock u2.mem\[128\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08727__I0 _03926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12502__CLK clknet_leaf_106_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07710_ u2.mem\[43\]\[10\] _03049_ _03050_ u2.mem\[20\]\[10\] _03179_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08690_ _03930_ u2.mem\[13\]\[11\] _03924_ _03931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_1456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08378__S _03733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10534__I0 _05018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07641_ _02502_ _03111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06902__A2 _02380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07572_ _02499_ _03043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09311_ _04327_ _00445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12652__CLK clknet_leaf_205_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06523_ _01988_ _02008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11532__S _05709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09242_ _04286_ _00417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06454_ _01913_ _01949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09173_ _04161_ u2.mem\[24\]\[10\] _04236_ _04239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13008__CLK clknet_leaf_240_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06385_ _01883_ _01884_ _01885_ _01886_ _01887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_120_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08124_ _03515_ _03561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11411__A1 _04071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08841__S _04024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11262__I1 u2.mem\[153\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08055_ _03510_ _03511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09736__I data_in_trans\[9\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07006_ _02483_ _02438_ _02439_ _02484_ _02485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__12032__CLK clknet_leaf_302_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11714__A2 _05808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07394__A2 _02866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09672__S _04549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06160__I _01666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08957_ _04096_ _04097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_103_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12182__CLK clknet_leaf_77_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08718__I0 _03917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07908_ _01973_ _03246_ _03352_ _03373_ _01490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_5_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08888_ _04050_ _04056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10525__I0 _05009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07146__A2 _02622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07839_ _02586_ _03306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10850_ _05282_ _01029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09143__I0 _04174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09509_ _04371_ u2.mem\[32\]\[6\] _04448_ _04451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10781_ _05241_ _01001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09694__I1 u2.mem\[36\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11442__S _05655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12520_ _00399_ clknet_leaf_118_clock u2.mem\[24\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12451_ _00330_ clknet_leaf_84_clock u2.mem\[20\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09446__I1 u2.mem\[30\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_244_clock_I clknet_5_19_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11402_ _05510_ _05631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06409__A1 _01878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12382_ _00261_ clknet_leaf_207_clock u2.mem\[16\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_165_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11333_ _05587_ u2.mem\[158\]\[1\] _05585_ _05588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11264_ _05499_ _05544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13003_ _00882_ clknet_leaf_249_clock u2.mem\[55\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12525__CLK clknet_leaf_188_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10215_ _04889_ u2.mem\[49\]\[1\] _04887_ _04890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11195_ _03491_ _05499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10146_ _04848_ _00759_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08709__I0 _03908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10521__S _05078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10077_ _04806_ u2.mem\[45\]\[10\] _04802_ _04807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08198__S _03609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10516__I0 _04998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09381__I _04147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07137__A2 _02371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09382__I0 _04371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09134__I0 _04161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10979_ _05366_ _01074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09685__I1 u2.mem\[36\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06648__A1 _01992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12718_ _00597_ clknet_leaf_252_clock u2.mem\[37\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12649_ _00528_ clknet_leaf_111_clock u2.mem\[32\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09437__I1 u2.mem\[30\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12055__CLK clknet_2_2__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11244__I1 u2.mem\[152\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06170_ _01608_ _01677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08661__S _03906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07073__A1 _02440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06820__A1 u2.mem\[144\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08948__I0 _04044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09860_ _04592_ u2.mem\[40\]\[8\] _04671_ _04672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13450__CLK clknet_leaf_343_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10755__I0 _05225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06179__A3 _01587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08811_ _03930_ u2.mem\[16\]\[11\] _04000_ _04004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09791_ _04602_ u2.mem\[38\]\[11\] _04628_ _04632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08742_ _03605_ _03606_ _03607_ _03878_ _03962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07128__A2 _02467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08176__I1 u2.mem\[2\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08673_ _03684_ _03919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10132__A1 _04417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06336__B1 _01680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_193_clock_I clknet_5_31_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07624_ _02623_ _03095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_311_clock clknet_5_17_0_clock clknet_leaf_311_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_53_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09125__I0 _04148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07555_ _02460_ _03026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11262__S _05536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06639__A1 u2.mem\[185\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06506_ _01990_ _01991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06639__B2 u2.mem\[173\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07486_ u2.mem\[23\]\[6\] _02913_ _02914_ u2.mem\[22\]\[6\] _02959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07300__A2 _02612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09225_ _04274_ u2.mem\[25\]\[10\] _04270_ _04275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06437_ _01769_ _01915_ _01932_ _01935_ _01466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_326_clock clknet_5_7_0_clock clknet_leaf_326_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09428__I1 u2.mem\[30\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09667__S _04544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09156_ _04229_ _00388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06368_ u2.mem\[191\]\[4\] _01681_ _01683_ u2.mem\[179\]\[4\] _01871_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08107_ _03549_ _00019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12548__CLK clknet_leaf_98_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07064__A1 u2.mem\[37\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09087_ _04189_ _00359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10606__S _05131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06299_ _01801_ _01802_ _01803_ _01804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_162_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10994__I0 _05340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08038_ _03497_ _03494_ _03498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06811__B2 u2.mem\[156\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08939__I0 _04035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11699__A1 _04120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10000_ _04714_ u2.mem\[43\]\[14\] _04755_ _04758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12698__CLK clknet_leaf_110_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09989_ _04703_ u2.mem\[43\]\[9\] _04750_ _04752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10341__S _04966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06327__B1 _01709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11951_ _05970_ _05971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11171__I0 _05464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06878__A1 _02347_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10902_ _05315_ _01048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11882_ _05928_ _05932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_3789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08746__S _03963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09116__I0 _04132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10833_ u2.mem\[63\]\[14\] _03533_ _05268_ _05271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12078__CLK clknet_leaf_343_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08545__I _03835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13552_ _01431_ clknet_leaf_13_clock u2.mem\[193\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10764_ _05231_ _05232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_164_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13323__CLK clknet_leaf_303_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12503_ _00382_ clknet_leaf_121_clock u2.mem\[23\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13483_ _01362_ clknet_leaf_290_clock u2.mem\[184\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09419__I1 u2.mem\[30\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10695_ _05115_ u2.mem\[60\]\[9\] _05184_ _05186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12434_ _00313_ clknet_leaf_124_clock u2.mem\[19\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12365_ _00244_ clknet_leaf_210_clock u2.mem\[15\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13473__CLK clknet_leaf_292_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10516__S _05073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11316_ _05577_ _01200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06802__A1 u2.mem\[188\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08280__I _03659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06802__B2 u2.mem\[187\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12296_ _00175_ clknet_leaf_120_clock u2.mem\[10\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11247_ _05534_ _01174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11178_ _05489_ _01150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10129_ _04838_ _00752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07624__I _02623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08158__I1 u2.mem\[2\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06318__B1 _01732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11162__I0 _05470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11146__I _05348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07530__A2 _02913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07340_ u2.mem\[49\]\[4\] _02660_ _02661_ u2.mem\[46\]\[4\] _02815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_91_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08455__I _03777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07271_ _02742_ _02743_ _02744_ _02746_ _02747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_91_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09010_ _04131_ _04132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06222_ _01565_ _01728_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07046__A1 _02466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06153_ _01570_ _01616_ _01644_ _01660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_145_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07597__A2 _03066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06084_ _01570_ _01591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12840__CLK clknet_leaf_139_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09912_ _04705_ u2.mem\[41\]\[10\] _04701_ _04706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09843_ _04662_ _00642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10161__S _04856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12990__CLK clknet_leaf_258_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06986_ _02464_ _02465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09774_ _04622_ _00613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09950__S _04729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08725_ _03923_ u2.mem\[14\]\[8\] _03952_ _03953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_250_clock clknet_5_22_0_clock clknet_leaf_250_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_2_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08656_ _03907_ _00210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12220__CLK clknet_leaf_215_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13346__CLK clknet_leaf_5_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07607_ _02592_ _03078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08587_ _03813_ u2.mem\[11\]\[6\] _03862_ _03865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07538_ u2.mem\[6\]\[7\] _02861_ _02862_ u2.mem\[47\]\[7\] _03010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_265_clock clknet_5_23_0_clock clknet_leaf_265_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_74_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07285__A1 u2.mem\[37\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07469_ _02938_ _02939_ _02940_ _02941_ _02942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__12370__CLK clknet_leaf_150_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13496__CLK clknet_leaf_312_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09208_ _04144_ _04263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10480_ _05050_ _05056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_108_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09139_ _04167_ u2.mem\[23\]\[12\] _04218_ _04219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07037__A1 _02407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10967__I0 _05343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08785__A1 _03983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12150_ _00029_ clknet_leaf_73_clock u2.mem\[1\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11101_ _05441_ _01121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12081_ net45 clknet_leaf_362_clock output_active_hold\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_203_clock clknet_5_29_0_clock clknet_leaf_203_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_104_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10719__I0 _05200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11032_ _05388_ u2.mem\[139\]\[3\] _05395_ _05399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06012__A2 _01517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10071__S _04802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_9_clock clknet_5_1_0_clock clknet_leaf_9_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_4232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09860__S _04671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_218_clock clknet_5_28_0_clock clknet_leaf_218_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_64_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11144__I0 _05468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12983_ _00862_ clknet_leaf_326_clock u2.mem\[53\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08476__S _03793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11934_ _05961_ _01434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11695__I1 u2.mem\[180\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11865_ _05909_ u2.mem\[191\]\[2\] _05918_ _05921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12713__CLK clknet_leaf_50_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08275__I _03491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10816_ _05261_ _01016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11796_ _04310_ _05847_ _05878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_43_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13535_ _01414_ clknet_leaf_329_clock u2.mem\[192\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10747_ _03704_ _05220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11630__S _05771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13466_ _01345_ clknet_leaf_347_clock u2.mem\[181\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10678_ _05176_ _00963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12863__CLK clknet_leaf_148_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_141_clock_I clknet_5_13_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07028__A1 _02441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12417_ _00296_ clknet_leaf_161_clock u2.mem\[18\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13397_ _01276_ clknet_leaf_307_clock u2.mem\[169\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12348_ _00227_ clknet_leaf_202_clock u2.mem\[14\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07043__A4 _02493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06787__B1 _02122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13219__CLK clknet_leaf_283_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12279_ _00158_ clknet_leaf_120_clock u2.mem\[9\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09576__I0 _04494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11383__I0 _05589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11077__S _05422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06679__B _02163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07200__A1 u2.mem\[28\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06840_ u2.mem\[165\]\[5\] _02075_ _02078_ u2.mem\[163\]\[5\] _02092_ u2.mem\[177\]\[5\]
+ _02320_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__06003__A2 _01510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07200__B2 u2.mem\[31\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12243__CLK clknet_leaf_73_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07354__I _02555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07751__A2 _03120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13369__CLK clknet_leaf_356_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06771_ u2.mem\[171\]\[3\] _02065_ _02067_ u2.mem\[157\]\[3\] _02253_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11135__I0 _05460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08510_ _03799_ _03818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_76_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09490_ _04438_ _00513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_66_clock_I clknet_5_3_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08441_ _03773_ _00129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06857__A4 _02336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06711__C2 u2.mem\[162\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08372_ _03732_ _00101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11438__I1 u2.mem\[164\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09500__I0 _04362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07323_ _02474_ _02798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07254_ u2.mem\[5\]\[2\] _02687_ _02688_ u2.mem\[38\]\[2\] _02731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07282__A4 _02757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07019__A1 _02410_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06205_ _01557_ _01586_ _01712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07185_ u2.mem\[43\]\[1\] _02515_ _02517_ u2.mem\[20\]\[1\] _02663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10156__S _04851_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06490__A2 _01933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06136_ _01642_ _01643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06242__A2 _01610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06067_ col_select_trans\[1\].data_sync _01574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_160_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09744__I data_in_trans\[11\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_343_clock_I clknet_5_5_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09826_ _04599_ u2.mem\[39\]\[10\] _04649_ _04652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09319__I0 _04285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07742__A2 _03031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09757_ data_in_trans\[14\].data_sync _04611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06969_ _02447_ _02448_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11126__I0 _05428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08708_ _03943_ _00226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08296__S _03660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09688_ _04491_ u2.mem\[36\]\[12\] _04559_ _04560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08639_ _03879_ _03895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11650_ _05662_ _05786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08095__I _03492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12886__CLK clknet_leaf_63_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10601_ _05132_ _00930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11581_ _05743_ _01299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11450__S _05654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10532_ _05016_ u2.mem\[56\]\[10\] _05083_ _05086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13320_ _01199_ clknet_leaf_306_clock u2.mem\[156\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08823__I _03987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12116__CLK clknet_leaf_328_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13251_ _01130_ clknet_leaf_285_clock u2.mem\[145\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10463_ _05046_ _00878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07439__I _02595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09855__S _04666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12202_ _00081_ clknet_leaf_54_clock u2.mem\[4\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13182_ _01061_ clknet_leaf_271_clock u2.mem\[133\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11601__I1 u2.mem\[174\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10394_ _04988_ _05002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_163_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07025__A4 _02434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12133_ _01459_ clknet_leaf_14_clock u2.driver_mem\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12266__CLK clknet_leaf_55_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12064_ data_in_trans\[7\].A clknet_leaf_300_clock data_in_trans\[7\].data_sync vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13511__CLK clknet_leaf_317_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11365__I0 _05583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11015_ _05345_ _05388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_157_clock clknet_5_26_0_clock clknet_leaf_157_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09590__S _04501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07733__A2 _03191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07107__C _02473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12966_ _00845_ clknet_leaf_87_clock u2.mem\[52\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08533__I1 u2.mem\[9\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07497__A1 _01945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11917_ _05907_ u2.mem\[193\]\[1\] _05950_ _05952_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12897_ _00776_ clknet_leaf_224_clock u2.mem\[48\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07123__B _02484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11848_ _05909_ u2.mem\[190\]\[2\] _05905_ _05910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11779_ _05864_ u2.mem\[186\]\[0\] _05866_ _05867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08733__I _03941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13518_ _01397_ clknet_leaf_330_clock u2.mem\[189\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_292_clock_I clknet_5_20_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13449_ _01328_ clknet_leaf_343_clock u2.mem\[178\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13041__CLK clknet_leaf_321_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12609__CLK clknet_leaf_155_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08990_ _04115_ _00336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07972__A2 _03425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13191__CLK clknet_leaf_279_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07941_ u2.mem\[17\]\[14\] _03310_ _03311_ u2.mem\[24\]\[14\] _03406_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12759__CLK clknet_leaf_50_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07872_ u2.mem\[1\]\[13\] _03261_ _03262_ u2.mem\[7\]\[13\] _03338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07185__B1 _02517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07724__A2 _03077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09611_ _04515_ _00557_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06823_ _02285_ _02290_ _02303_ _02304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_83_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11108__I0 _05424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11535__S _05709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09542_ _04135_ _04471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06754_ u2.mem\[169\]\[2\] _02141_ _02143_ u2.mem\[147\]\[2\] _02236_ _02237_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__11659__I1 u2.mem\[178\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08524__I1 u2.mem\[9\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09721__I0 _04583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09473_ _04418_ _04429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07488__B2 u2.mem\[21\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06685_ _02167_ _02168_ _02169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08424_ _03753_ _03764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_145_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08844__S _04024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06428__I _01927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12139__CLK clknet_leaf_212_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08355_ _03720_ _00096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11270__S _05546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07306_ u2.mem\[45\]\[4\] _02633_ _02634_ u2.mem\[34\]\[4\] _02781_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08286_ _03664_ u2.mem\[5\]\[1\] _03660_ _03665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11831__I1 u2.mem\[189\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06999__B1 _02477_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07237_ _02710_ _02711_ _02712_ _02713_ _02714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_137_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06463__A2 _01931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12289__CLK clknet_leaf_165_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07168_ _02504_ _02646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13534__CLK clknet_leaf_318_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11595__I0 _05752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07412__A1 _02880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06119_ u2.mem\[184\]\[0\] _01625_ _01553_ _01626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08460__I0 _03685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07099_ _02419_ _02578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_78_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_74_clock clknet_5_8_0_clock clknet_leaf_74_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07963__A2 _02509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11898__I1 _03521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09809_ _04642_ _00628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_89_clock clknet_5_10_0_clock clknet_leaf_89_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12820_ _00699_ clknet_leaf_61_clock u2.mem\[43\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09712__I0 _04576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12751_ _00630_ clknet_leaf_225_clock u2.mem\[39\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11702_ _05819_ _01344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_12_clock clknet_5_3_0_clock clknet_leaf_12_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12682_ _00561_ clknet_leaf_127_clock u2.mem\[34\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11633_ _05776_ _01318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09649__I _04521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11564_ _05713_ u2.mem\[172\]\[2\] _05731_ _05734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_27_clock clknet_5_2_0_clock clknet_leaf_27_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_11_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13303_ _01182_ clknet_leaf_362_clock u2.mem\[154\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10515_ _05076_ _00900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11495_ _04223_ _05690_ _05691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_171_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_14_clock_I clknet_5_3_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13234_ _01113_ clknet_leaf_278_clock u2.mem\[142\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10446_ _05005_ u2.mem\[54\]\[5\] _05035_ _05037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08451__I0 _03668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13165_ _01044_ clknet_leaf_264_clock u2.mem\[131\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10377_ _04988_ _04989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12901__CLK clknet_leaf_74_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09384__I _04150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12116_ _01479_ clknet_leaf_328_clock u2.select_mem_row\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13096_ _00975_ clknet_leaf_47_clock u2.mem\[60\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12047_ net6 clknet_2_2__leaf_clock_a col_select_trans\[5\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07118__B _02507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11889__I1 _03511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_239_clock_I clknet_5_19_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11355__S _05598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06390__B2 u2.mem\[188\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12949_ _00828_ clknet_leaf_67_clock u2.mem\[51\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13407__CLK clknet_leaf_304_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06470_ _01958_ _01955_ _01959_ _01961_ _01473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_61_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08664__S _03906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06142__A1 _01612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07485__A4 _02957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11090__S _05435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10077__I0 _04806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09559__I _04464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08140_ _03528_ _03572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11813__I1 u2.mem\[188\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06445__A2 _01931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08071_ _01958_ _03517_ _03522_ _00010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08690__I0 _03930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07022_ u2.mem\[58\]\[0\] _02495_ _02500_ u2.mem\[36\]\[0\] _02501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12581__CLK clknet_leaf_98_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09294__I _04312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07945__A2 _02627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08973_ _04030_ u2.mem\[20\]\[7\] _04102_ _04106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11329__I _05584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10233__I _04588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07924_ u2.mem\[44\]\[14\] _02521_ _02523_ u2.mem\[42\]\[14\] _03389_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07855_ _02618_ _03322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06806_ u2.mem\[180\]\[4\] _02043_ _02014_ u2.mem\[172\]\[4\] _02287_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07786_ u2.mem\[40\]\[12\] _03251_ _03252_ u2.mem\[30\]\[12\] _03253_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07542__I _02360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06381__B2 u2.mem\[164\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09525_ _04387_ u2.mem\[32\]\[13\] _04458_ _04460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06737_ u2.mem\[165\]\[2\] _02076_ _02079_ u2.mem\[163\]\[2\] u2.mem\[145\]\[2\]
+ _02081_ _02220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_37_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11501__I0 _05671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13087__CLK clknet_leaf_245_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08574__S _03857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09456_ _04356_ u2.mem\[31\]\[0\] _04419_ _04420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06668_ _02152_ _02153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07330__B1 _02649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_08407_ _03657_ u2.mem\[7\]\[0\] _03754_ _03755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09387_ _04153_ _04375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06599_ _02023_ _02058_ _02084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08373__I _03727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08338_ _03706_ u2.mem\[5\]\[11\] _03694_ _03707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11804__I1 u2.mem\[187\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08269_ _03575_ u2.mem\[4\]\[13\] _03650_ _03652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10408__I _04988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07633__B2 u2.mem\[30\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08681__I0 _03923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12924__CLK clknet_leaf_257_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10300_ _04943_ _04944_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_leaf_188_clock_I clknet_5_31_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11280_ _05555_ _01186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06841__C1 u2.mem\[193\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11568__I0 _05717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10231_ _04900_ u2.mem\[49\]\[6\] _04896_ _04901_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10162_ _04857_ _00766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10093_ _04817_ u2.mem\[45\]\[15\] _04811_ _04818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_240_clock_I clknet_5_19_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08736__I1 u2.mem\[14\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12304__CLK clknet_leaf_164_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11175__S _05484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06372__A1 _01867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12803_ _00682_ clknet_leaf_145_clock u2.mem\[42\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10995_ _05375_ _01081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11903__S _05942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12010__D mem_address_trans\[2\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12734_ _00613_ clknet_leaf_252_clock u2.mem\[38\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12454__CLK clknet_leaf_85_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06675__A2 _02154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12665_ _00544_ clknet_leaf_58_clock u2.mem\[33\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10519__S _05078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11616_ _05756_ u2.mem\[175\]\[4\] _05760_ _05766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08283__I _03496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12596_ _00475_ clknet_leaf_99_clock u2.mem\[29\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10318__I _04943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11547_ _05711_ u2.mem\[171\]\[1\] _05722_ _05724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11478_ _05680_ u2.mem\[166\]\[5\] _05664_ _05681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13217_ _01096_ clknet_leaf_286_clock u2.mem\[139\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10429_ _05026_ _00864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10231__I0 _04900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13148_ _01027_ clknet_leaf_263_clock u2.mem\[128\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11149__I _05351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13079_ _00958_ clknet_leaf_43_clock u2.mem\[59\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08727__I1 u2.mem\[14\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11731__I0 _05837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07640_ _03106_ _03107_ _03108_ _03109_ _03110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_54_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07362__I _02581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07571_ _02494_ _03042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09310_ _04276_ u2.mem\[27\]\[11\] _04323_ _04327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06522_ _02006_ _02007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11813__S _05888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06115__A1 _01571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09241_ _04285_ u2.mem\[25\]\[15\] _04279_ _04286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06453_ _01918_ _01948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12947__CLK clknet_leaf_233_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09172_ _04238_ _00395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08193__I mem_address_trans\[1\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06384_ u2.mem\[184\]\[5\] _01778_ _01749_ _01886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11798__I0 _05864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08123_ _03560_ _00024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07615__A1 _03076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11411__A2 _05606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08054_ data_in_trans\[5\].data_sync _03510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07005_ _02440_ _02441_ _02382_ _02484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_134_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07379__B1 _02688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06441__I _01914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12327__CLK clknet_leaf_126_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08956_ _04095_ _03988_ _04096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_88_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input30_I mem_address_a[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09915__I0 _04707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07907_ _03357_ _03362_ _03367_ _03372_ _03373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_3905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08887_ _04055_ _00293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11722__I0 _05831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07838_ _02584_ _03305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06354__A1 u2.mem\[187\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12477__CLK clknet_leaf_181_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06354__B2 u2.mem\[192\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07769_ u2.mem\[52\]\[11\] _03080_ _03081_ u2.mem\[21\]\[11\] _03237_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09508_ _04450_ _00519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10780_ _05211_ u2.mem\[62\]\[7\] _05237_ _05241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_09439_ _04380_ u2.mem\[30\]\[10\] _04406_ _04409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10339__S _04966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_12450_ _00329_ clknet_leaf_159_clock u2.mem\[20\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11401_ _05630_ _01232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06409__A2 _01554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12381_ _00260_ clknet_leaf_206_clock u2.mem\[16\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_165_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11332_ _05504_ _05587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10074__S _04802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11263_ _05543_ _01181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07909__A2 _02444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13002_ _00881_ clknet_leaf_322_clock u2.mem\[54\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10214_ _04569_ _04889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11194_ _05498_ _01157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10145_ _04795_ u2.mem\[47\]\[5\] _04846_ _04848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12005__D net24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13252__CLK clknet_leaf_291_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10802__S _05253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06593__A1 _02031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08709__I1 u2.mem\[14\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09906__I0 _04700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10076_ _04598_ _04806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10516__I1 u2.mem\[56\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08278__I _03541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07182__I _02530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_10978_ _05335_ u2.mem\[136\]\[0\] _05365_ _05366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06648__A2 _02052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12717_ _00596_ clknet_leaf_254_clock u2.mem\[37\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08893__I0 _04028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12648_ _00527_ clknet_leaf_114_clock u2.mem\[32\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12579_ _00458_ clknet_leaf_104_clock u2.mem\[28\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06281__B1 _01631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09773__S _04618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08810_ _04003_ _00268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11808__S _05878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08389__S _03738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09790_ _04631_ _00620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06584__A1 u2.mem\[171\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09572__I _04464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06584__B2 u2.mem\[157\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08741_ _03961_ _00241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11607__I _05760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08672_ _03918_ _00215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_136_clock_I clknet_5_13_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06336__A1 u2.mem\[147\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10132__A2 _04760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07623_ _02621_ _03094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07554_ _02456_ _03025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08916__I _04071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06505_ _01988_ _01989_ _01990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07485_ _02954_ _02955_ _02956_ _02957_ _02958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_107_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08884__I0 _04019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09224_ _04160_ _04274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06436_ u2.mem\[193\]\[2\] _01928_ _01933_ u2.mem\[194\]\[2\] _01934_ _01935_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_22_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13125__CLK clknet_leaf_23_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09155_ _04132_ u2.mem\[24\]\[2\] _04226_ _04229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06367_ u2.mem\[170\]\[4\] _01686_ _01688_ u2.mem\[156\]\[4\] _01870_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08106_ _03548_ u2.mem\[1\]\[1\] _03546_ _03549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07064__A2 _02540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09086_ _04145_ u2.mem\[22\]\[5\] _04187_ _04189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06298_ u2.mem\[146\]\[2\] _01692_ _01694_ u2.mem\[186\]\[2\] _01803_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08037_ _03496_ _03497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_150_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09683__S _04554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06171__I _01677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09061__I0 _04171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11699__A2 _05808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10622__S _05141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09988_ _04751_ _00698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09482__I _04418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07772__B1 _03154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08939_ _04035_ u2.mem\[19\]\[9\] _04084_ _04086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10421__I _04988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08098__I _03541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11950_ _03582_ _05926_ _05970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06327__A1 u2.mem\[153\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06327__B2 u2.mem\[160\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11171__I1 u2.mem\[148\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10901_ _05305_ u2.mem\[131\]\[4\] _05309_ _05315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06878__A2 _02351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11881_ _05931_ _01411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10832_ _05270_ _01023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13551_ _01430_ clknet_leaf_13_clock u2.mem\[193\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10763_ _04394_ _05172_ _05231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_12502_ _00381_ clknet_leaf_106_clock u2.mem\[23\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_338_clock_I clknet_5_5_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08762__S _03973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13482_ _01361_ clknet_leaf_298_clock u2.mem\[183\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10694_ _05185_ _00970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12433_ _00312_ clknet_leaf_161_clock u2.mem\[19\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07055__A2 _02531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12364_ _00243_ clknet_leaf_206_clock u2.mem\[15\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11315_ _05544_ u2.mem\[157\]\[0\] _05576_ _05577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12295_ _00174_ clknet_leaf_120_clock u2.mem\[10\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06081__I _01587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09052__I0 _04164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11246_ _05514_ u2.mem\[152\]\[4\] _05528_ _05534_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11628__S _05771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10532__S _05083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11177_ _05470_ u2.mem\[148\]\[4\] _05483_ _05489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07763__B1 _03067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10128_ _04815_ u2.mem\[46\]\[14\] _04835_ _04838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11427__I _05646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12792__CLK clknet_leaf_44_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10059_ _04794_ _00726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07126__B _02393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06318__A1 u2.mem\[145\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08937__S _04084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07515__B1 _02891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06318__B2 u2.mem\[168\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11162__I1 u2.mem\[147\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12022__CLK clknet_leaf_287_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13148__CLK clknet_leaf_263_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07270_ u2.mem\[3\]\[3\] _02480_ _02745_ _02746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_149_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07294__A2 _02591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06221_ _01726_ _01727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12172__CLK clknet_leaf_210_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10425__I0 _05023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06152_ _01658_ _01659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07046__A2 _02467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_62_clock_I clknet_5_9_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06254__B1 _01666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06083_ u2.mem\[177\]\[0\] _01583_ _01589_ u2.mem\[168\]\[0\] _01590_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07087__I _02417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09911_ _04598_ _04705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11538__S _05708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09842_ _04565_ u2.mem\[40\]\[0\] _04661_ _04662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06557__A1 _02041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07754__B1 _03050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07815__I _02514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09773_ _04576_ u2.mem\[38\]\[3\] _04618_ _04622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_06985_ _02458_ _02459_ _02463_ _02398_ _02464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08724_ _03941_ _03952_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_85_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06309__A1 u2.mem\[184\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_287_clock_I clknet_5_20_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08847__S _04024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_14_0_clock clknet_3_7_0_clock clknet_4_14_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_54_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08655_ _03900_ u2.mem\[13\]\[0\] _03906_ _03907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11273__S _05546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07606_ _02590_ _03077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06324__A4 _01827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08586_ _03864_ _00183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07550__I _02427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07537_ u2.mem\[8\]\[7\] _02858_ _02859_ u2.mem\[4\]\[7\] _03009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08857__I0 _04035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12515__CLK clknet_leaf_105_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10664__I0 _05121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06166__I _01672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07468_ u2.mem\[58\]\[6\] _02809_ _02810_ u2.mem\[36\]\[6\] _02941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07285__A2 _02540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09207_ _04262_ _00406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06419_ _01913_ _01920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07399_ u2.mem\[15\]\[5\] _02792_ _02793_ u2.mem\[13\]\[5\] _02873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09138_ _04202_ _04218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07037__A2 _02408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12665__CLK clknet_leaf_58_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09069_ _04177_ u2.mem\[21\]\[15\] _04168_ _04178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11100_ _05432_ u2.mem\[143\]\[5\] _05434_ _05441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12080_ data_in_trans\[15\].A clknet_leaf_303_clock data_in_trans\[15\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06260__A3 _01765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10719__I1 u2.mem\[61\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11448__S _05655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11031_ _05398_ _01094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10151__I _04840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08757__S _03968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12045__CLK clknet_2_2__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12982_ _00861_ clknet_leaf_31_clock u2.mem\[53\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09940__I _04718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11144__I1 u2.mem\[146\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11933_ _05213_ u2.mem\[193\]\[8\] _05960_ _05961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11183__S _05492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11864_ _05920_ _01405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06720__A1 _02179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12195__CLK clknet_leaf_72_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10815_ u2.mem\[63\]\[6\] _03513_ _05258_ _05261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11795_ _05877_ _01379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09588__S _04501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10655__I0 _05112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13440__CLK clknet_leaf_341_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13534_ _01413_ clknet_leaf_318_clock u2.mem\[192\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10746_ _05219_ _00988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13465_ _01344_ clknet_leaf_346_clock u2.mem\[181\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10677_ _05097_ u2.mem\[60\]\[1\] _05174_ _05176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09387__I _04153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12416_ _00295_ clknet_leaf_160_clock u2.mem\[18\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07028__A2 _02382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13396_ _01275_ clknet_leaf_310_clock u2.mem\[169\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11080__I0 _05428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12347_ _00226_ clknet_leaf_221_clock u2.mem\[14\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06787__A1 u2.mem\[146\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06787__B2 u2.mem\[173\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_310_clock clknet_5_17_0_clock clknet_leaf_310_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12278_ _00157_ clknet_leaf_101_clock u2.mem\[9\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11229_ _05511_ u2.mem\[151\]\[3\] _05520_ _05524_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11383__I1 u2.mem\[161\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07200__A2 _02585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_325_clock clknet_5_7_0_clock clknet_leaf_325_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_7_1462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06770_ u2.mem\[167\]\[3\] _02060_ _02062_ u2.mem\[183\]\[3\] _02252_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09850__I _04660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11135__I1 u2.mem\[146\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12538__CLK clknet_leaf_115_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08440_ _03723_ u2.mem\[7\]\[15\] _03769_ _03773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06711__A1 u2.mem\[154\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07370__I _02592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06711__B2 u2.mem\[148\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08371_ _03672_ u2.mem\[6\]\[3\] _03728_ _03732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11821__S _05887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09500__I1 u2.mem\[32\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07322_ u2.mem\[1\]\[4\] _02795_ _02796_ u2.mem\[7\]\[4\] _02797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10646__I0 _05103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07253_ _02726_ _02727_ _02728_ _02729_ _02730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_104_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10437__S _05030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06204_ u2.mem\[153\]\[0\] _01708_ _01710_ u2.mem\[160\]\[0\] _01711_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07184_ u2.mem\[49\]\[1\] _02660_ _02661_ u2.mem\[46\]\[1\] _02662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07019__A2 _02391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06714__I _02133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11071__I0 _05420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06227__B1 _01732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06135_ _01641_ _01596_ _01642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09016__I0 _04136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06066_ col_select_trans\[0\].data_sync _01573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12068__CLK clknet_leaf_33_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07545__I _02395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09961__S _04734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09825_ _04651_ _00635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13313__CLK clknet_leaf_349_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09756_ _04610_ _00607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06968_ _02429_ _02445_ _02446_ _02393_ _02447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__11126__I1 u2.mem\[145\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08707_ _03900_ u2.mem\[14\]\[0\] _03942_ _03943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09687_ _04543_ _04559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_2_1__f_clock_a clknet_0_clock_a clknet_2_1__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_27_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06899_ _02377_ _02378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_2127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13463__CLK clknet_leaf_344_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08638_ _03894_ _00205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08569_ _03854_ _00176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10637__I0 _05093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10600_ _05093_ u2.mem\[58\]\[0\] _05131_ _05132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11580_ _05715_ u2.mem\[173\]\[3\] _05739_ _05743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10262__A1 _03583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10531_ _05085_ _00907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13250_ _01129_ clknet_leaf_285_clock u2.mem\[145\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10462_ _05020_ u2.mem\[54\]\[12\] _05045_ _05046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09000__I _04123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12201_ _00080_ clknet_leaf_54_clock u2.mem\[4\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11062__I0 _05388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13181_ _01060_ clknet_leaf_271_clock u2.mem\[133\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06769__A1 u2.mem\[164\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10393_ _05000_ _05001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11762__A1 _04248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06769__B2 u2.mem\[178\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12132_ _01473_ clknet_leaf_34_clock u2.driver_mem\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12063_ net20 clknet_2_3__leaf_clock_a data_in_trans\[7\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07718__B1 _03140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11365__I1 u2.mem\[160\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11014_ _05387_ _01088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07194__A1 _02668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07733__A3 _03196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_10_clock_I clknet_5_1_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12965_ _00844_ clknet_leaf_85_clock u2.mem\[52\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11916_ _05951_ _01426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12896_ _00775_ clknet_leaf_224_clock u2.mem\[48\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12830__CLK clknet_leaf_220_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07123__C _02483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11847_ _03666_ _05909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07249__A2 _02680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11778_ _05865_ _05866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_53_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13517_ _01396_ clknet_leaf_318_clock u2.mem\[189\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10729_ _05207_ u2.mem\[61\]\[5\] _05205_ _05208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_235_clock_I clknet_5_18_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12980__CLK clknet_leaf_43_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13448_ _01327_ clknet_leaf_343_clock u2.mem\[178\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08950__S _04089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10005__A1 _04334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06209__B1 _01715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13379_ _01258_ clknet_leaf_352_clock u2.mem\[166\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12210__CLK clknet_leaf_232_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13336__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07421__A2 _02893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07940_ u2.mem\[23\]\[14\] _02596_ _02598_ u2.mem\[22\]\[14\] _03405_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07972__A3 _03430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07709__B1 _03127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07365__I _02586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_264_clock clknet_5_23_0_clock clknet_leaf_264_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_155_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07871_ u2.mem\[15\]\[13\] _03258_ _03259_ u2.mem\[13\]\[13\] _03337_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_151_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07185__B2 u2.mem\[20\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09610_ _04489_ u2.mem\[34\]\[11\] _04511_ _04515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12360__CLK clknet_leaf_136_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13486__CLK clknet_leaf_298_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06822_ _02295_ _02300_ _02301_ _02302_ _02303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_68_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06932__A1 _02410_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11108__I1 u2.mem\[144\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09541_ _04470_ _00532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06753_ _02233_ _02234_ _02235_ _02236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_leaf_279_clock clknet_5_21_0_clock clknet_leaf_279_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_36_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09472_ _04428_ _00505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06684_ u2.mem\[179\]\[1\] _02151_ _02153_ u2.mem\[191\]\[1\] _02168_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08423_ _03763_ _00121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_202_clock clknet_5_29_0_clock clknet_leaf_202_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11551__S _05722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08354_ _03719_ u2.mem\[5\]\[14\] _03711_ _03720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09485__I0 _04387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07305_ _02360_ _02780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06448__B1 _01943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11292__I0 _05552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10167__S _04856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08285_ _03663_ _03664_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09956__S _04729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_8_clock clknet_5_1_0_clock clknet_leaf_8_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07236_ u2.mem\[43\]\[2\] _02515_ _02517_ u2.mem\[20\]\[2\] _02713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_153_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08860__S _04033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_217_clock clknet_5_28_0_clock clknet_leaf_217_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_164_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07167_ _02502_ _02645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_173_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06118_ _01586_ _01617_ _01625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_160_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07098_ _02417_ _02577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__08460__I1 u2.mem\[8\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12703__CLK clknet_leaf_239_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06049_ _01550_ _01551_ _01556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_132_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09808_ _04573_ u2.mem\[39\]\[2\] _04639_ _04642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12853__CLK clknet_leaf_80_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09739_ _04597_ _00603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_184_clock_I clknet_5_27_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11525__I _05708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10858__I0 _05194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12750_ _00629_ clknet_leaf_213_clock u2.mem\[39\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09712__I1 u2.mem\[37\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11701_ _05786_ u2.mem\[181\]\[0\] _05818_ _05819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12681_ _00560_ clknet_leaf_129_clock u2.mem\[34\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13209__CLK clknet_leaf_281_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06151__A2 _01609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11632_ _05756_ u2.mem\[176\]\[4\] _05770_ _05776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09476__I0 _04378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06439__B1 _01933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10077__S _04802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11563_ _05733_ _01291_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09866__S _04671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13302_ _01181_ clknet_leaf_7_clock u2.mem\[153\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10514_ _04995_ u2.mem\[56\]\[2\] _05073_ _05076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09228__I0 _04276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12233__CLK clknet_leaf_57_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13359__CLK clknet_leaf_357_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11494_ _05605_ _05690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_143_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13233_ _01112_ clknet_leaf_285_clock u2.mem\[142\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12008__D mem_address_trans\[1\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10445_ _05036_ _00870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13164_ _01043_ clknet_leaf_270_clock u2.mem\[130\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10376_ _04121_ _04964_ _04988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_87_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12383__CLK clknet_leaf_223_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12115_ _01478_ clknet_leaf_332_clock u2.select_mem_row\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13095_ _00974_ clknet_leaf_46_clock u2.mem\[60\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06303__B _01807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12046_ col_select_trans\[4\].A clknet_leaf_288_clock col_select_trans\[4\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07118__C _02426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07706__A3 _03173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09106__S _04197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06390__A2 _01601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07134__B _02498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10849__I0 _05202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12948_ _00827_ clknet_leaf_66_clock u2.mem\[51\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06529__I _02013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12879_ _00758_ clknet_leaf_230_clock u2.mem\[47\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09467__I0 _04369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09219__I0 _04269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06264__I _01768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08070_ _03521_ _03519_ _03522_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07021_ _02499_ _02500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11026__I0 _05380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06850__B1 _02122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12726__CLK clknet_leaf_72_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09575__I _04170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08972_ _04105_ _00328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12876__CLK clknet_leaf_215_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07923_ _03384_ _03385_ _03386_ _03387_ _03388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_116_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07158__A1 u2.mem\[32\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07158__B2 u2.mem\[2\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07854_ _02616_ _03321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10450__S _05035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09016__S _04124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06805_ u2.mem\[176\]\[4\] _02004_ _02020_ u2.mem\[189\]\[4\] _02286_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07785_ _02414_ _03252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12106__CLK clknet_leaf_58_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09524_ _04459_ _00526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06736_ u2.mem\[166\]\[2\] _02097_ _02099_ u2.mem\[161\]\[2\] _02218_ _02219_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_71_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_141_clock clknet_5_13_0_clock clknet_leaf_141_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09455_ _04418_ _04419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_06667_ _02104_ _01999_ _02152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_08406_ _03753_ _03754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_52_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08654__I _03905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09386_ _04374_ _00473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09458__I0 _04360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12256__CLK clknet_leaf_228_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07881__A2 _02521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06598_ u2.mem\[165\]\[0\] _02076_ _02079_ u2.mem\[163\]\[0\] u2.mem\[145\]\[0\]
+ _02082_ _02083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_24_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13501__CLK clknet_leaf_330_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08337_ _03705_ _03706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_156_clock clknet_5_26_0_clock clknet_leaf_156_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_123_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08268_ _03651_ _00078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07219_ u2.mem\[32\]\[2\] _02386_ _02396_ u2.mem\[2\]\[2\] _02696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06841__C2 _02089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08199_ _03610_ _00050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11568__I1 u2.mem\[172\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10230_ _04585_ _04900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07397__A1 u2.mem\[27\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10161_ _04810_ u2.mem\[47\]\[12\] _04856_ _04857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10424__I _03713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10092_ _04614_ _04817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06372__A2 _01868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13031__CLK clknet_leaf_326_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12802_ _00681_ clknet_leaf_145_clock u2.mem\[42\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10994_ _05340_ u2.mem\[137\]\[1\] _05373_ _05375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_109_clock clknet_5_11_0_clock clknet_leaf_109_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12733_ _00612_ clknet_leaf_255_clock u2.mem\[38\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12664_ _00543_ clknet_leaf_135_clock u2.mem\[33\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13181__CLK clknet_leaf_271_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11615_ _05765_ _01311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12595_ _00474_ clknet_leaf_105_clock u2.mem\[29\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12749__CLK clknet_leaf_212_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06084__I _01570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11546_ _05723_ _01284_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11477_ _05679_ _05680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_5_22_0_clock_I clknet_4_11_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13216_ _01095_ clknet_leaf_282_clock u2.mem\[139\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10428_ _05025_ u2.mem\[53\]\[14\] _05021_ _05026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12899__CLK clknet_leaf_64_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13147_ _01026_ clknet_leaf_265_clock u2.mem\[128\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10359_ _04907_ u2.mem\[52\]\[9\] _04976_ _04978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13078_ _00957_ clknet_leaf_25_clock u2.mem\[59\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12129__CLK clknet_leaf_35_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10270__S _04923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12029_ net39 clknet_2_2__leaf_clock_a row_select_trans\[2\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11731__I1 u2.mem\[182\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07570_ u2.mem\[53\]\[8\] _03039_ _03040_ u2.mem\[56\]\[8\] _03041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12279__CLK clknet_leaf_120_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09688__I0 _04491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06521_ _02005_ row_select_trans\[4\].data_sync _02006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13524__CLK clknet_leaf_15_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06115__A2 _01607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07312__B2 u2.mem\[30\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09240_ _04176_ _04285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06452_ u2.mem\[194\]\[6\] _01946_ _01947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07863__A2 _03323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_73_clock clknet_5_8_0_clock clknet_leaf_73_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_146_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09171_ _04158_ u2.mem\[24\]\[9\] _04236_ _04238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06383_ u2.mem\[171\]\[5\] _01610_ _01770_ u2.mem\[157\]\[5\] _01885_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10509__I _05072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08112__I0 _03552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08122_ _03559_ u2.mem\[1\]\[6\] _03555_ _03560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11798__I1 u2.mem\[187\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09860__I0 _04592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_132_clock_I clknet_5_12_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08053_ _01844_ _03505_ _03509_ _00005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_88_clock clknet_5_10_0_clock clknet_leaf_88_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07004_ _02412_ _02483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_162_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_11_clock clknet_5_3_0_clock clknet_leaf_11_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_66_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08955_ _04094_ _04095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_130_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11276__S _05546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13054__CLK clknet_leaf_259_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07906_ _03368_ _03369_ _03370_ _03371_ _03372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_44_1566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10180__S _04865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08886_ _04021_ u2.mem\[18\]\[3\] _04051_ _04055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input23_I inverter_select_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11722__I1 u2.mem\[182\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07837_ u2.mem\[9\]\[12\] _03302_ _03303_ u2.mem\[25\]\[12\] _03304_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_3928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_26_clock clknet_5_2_0_clock clknet_leaf_26_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06169__I _01675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07768_ u2.mem\[17\]\[11\] _03077_ _03078_ u2.mem\[24\]\[11\] _03236_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09679__I0 _04482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_57_clock_I clknet_5_12_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09507_ _04369_ u2.mem\[32\]\[5\] _04448_ _04450_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11486__I0 _05671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06719_ _02195_ _02197_ _02201_ _02202_ _02203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_38_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07699_ u2.mem\[16\]\[10\] _03031_ _03032_ u2.mem\[33\]\[10\] _03168_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07303__A1 _02763_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_09438_ _04408_ _00491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_09369_ _04362_ u2.mem\[29\]\[2\] _04358_ _04363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08103__I0 _03539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11400_ _05629_ u2.mem\[162\]\[2\] _05625_ _05630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12380_ _00259_ clknet_leaf_205_clock u2.mem\[16\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09851__I0 _04579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11331_ _05586_ _01206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06814__B1 _02144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06290__A1 u2.mem\[153\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11262_ _05517_ u2.mem\[153\]\[5\] _05536_ _05543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06290__B2 u2.mem\[160\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06632__I _02116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13001_ _00880_ clknet_leaf_322_clock u2.mem\[54\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10213_ _04888_ _00786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11193_ _05472_ u2.mem\[149\]\[5\] _05491_ _05498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10144_ _04847_ _00758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06593__A2 _02077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_334_clock_I clknet_5_6_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10075_ _04805_ _00731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07137__A4 _02468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13547__CLK clknet_leaf_35_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06345__A2 _01846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10977_ _05364_ _05365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_43_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12571__CLK clknet_leaf_182_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11713__I _03655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12716_ _00595_ clknet_leaf_254_clock u2.mem\[37\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08294__I _03670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12647_ _00526_ clknet_leaf_114_clock u2.mem\[32\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12578_ _00457_ clknet_leaf_169_clock u2.mem\[28\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09842__I0 _04565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11529_ _05711_ u2.mem\[170\]\[1\] _05709_ _05712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06281__B2 u2.mem\[188\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13077__CLK clknet_leaf_25_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07230__B1 _02489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11096__S _05435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06698__B _01993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08740_ _03939_ u2.mem\[14\]\[15\] _03957_ _03961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07373__I _02602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08671_ _03917_ u2.mem\[13\]\[5\] _03915_ _03918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06336__A2 _01676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07533__B2 u2.mem\[19\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07622_ u2.mem\[8\]\[8\] _03091_ _03092_ u2.mem\[4\]\[8\] _03093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12914__CLK clknet_leaf_157_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07553_ _03014_ _03017_ _03020_ _03023_ _03024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_81_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08333__I0 _03702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11623__I _05770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06504_ row_select_trans\[3\].data_sync _01989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07484_ u2.mem\[28\]\[6\] _02839_ _02840_ u2.mem\[31\]\[6\] _02957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10140__I0 _04790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09223_ _04273_ _00411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06435_ _01920_ _01934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09154_ _04228_ _00387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06366_ u2.mem\[173\]\[4\] _01719_ _01721_ u2.mem\[185\]\[4\] _01869_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09833__I0 _04609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_283_clock_I clknet_5_21_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_10_0_clock clknet_3_5_0_clock clknet_4_10_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08105_ _03497_ _03548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11640__I0 _05750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09085_ _04188_ _00358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06297_ u2.mem\[191\]\[2\] _01682_ _01684_ u2.mem\[179\]\[2\] _01802_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07548__I _02414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06272__A1 u2.mem\[167\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08036_ data_in_trans\[1\].data_sync _03496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06272__B2 u2.mem\[183\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09061__I1 u2.mem\[21\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10903__S _05309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06024__A1 u2.driver_mem\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07221__B1 _02436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12444__CLK clknet_leaf_198_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07367__A4 _02841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09987_ _04700_ u2.mem\[43\]\[8\] _04750_ _04751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07772__B2 u2.mem\[38\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08938_ _04085_ _00314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08869_ _03714_ _04044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06327__A2 _01707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10900_ _05314_ _01047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11880_ u2.mem\[192\]\[1\] _03497_ _05929_ _05931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06878__A3 _02356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10831_ u2.mem\[63\]\[13\] _03531_ _05268_ _05270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07288__B1 _02674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13550_ _01429_ clknet_leaf_12_clock u2.mem\[193\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10762_ _05230_ _00993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09003__I data_in_trans\[1\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12501_ _00380_ clknet_leaf_106_clock u2.mem\[23\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13481_ _01360_ clknet_leaf_296_clock u2.mem\[183\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10693_ _05112_ u2.mem\[60\]\[8\] _05184_ _05185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12432_ _00311_ clknet_leaf_159_clock u2.mem\[19\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09824__I0 _04596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12363_ _00242_ clknet_leaf_208_clock u2.mem\[15\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11314_ _05575_ _05576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_4_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12294_ _00173_ clknet_leaf_101_clock u2.mem\[10\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11909__S _05928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11245_ _05533_ _01173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12016__D mem_address_trans\[5\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10198__I0 _04808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06015__A1 u2.driver_mem\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07212__B1 _02619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11176_ _05488_ _01149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07763__A1 u2.mem\[29\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10127_ _04837_ _00751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12937__CLK clknet_leaf_323_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08289__I _03666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10058_ _04792_ u2.mem\[45\]\[4\] _04793_ _04794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07126__C _02547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07515__A1 u2.mem\[14\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07515__B2 u2.mem\[12\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11644__S _05779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10370__I0 _04918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09114__S _04203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07279__B1 _02661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07142__B _02507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12317__CLK clknet_leaf_197_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06981__B _02442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06220_ u2.mem\[0\]\[1\] _01726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08752__I _03962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09815__I0 _04583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06151_ _01567_ _01609_ _01658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10425__I1 u2.mem\[53\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06254__A1 u2.mem\[180\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12467__CLK clknet_leaf_108_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06254__B2 u2.mem\[150\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06082_ _01586_ _01588_ _01589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_171_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11819__S _05888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09910_ _04704_ _00667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10189__I0 _04799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09841_ _04660_ _04661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_113_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06557__A2 _02000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07754__B2 u2.mem\[20\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09772_ _04621_ _00612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06984_ _02440_ _02401_ _02382_ _02463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XTAP_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08723_ _03951_ _00233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11689__I0 _05790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08654_ _03905_ _03906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08927__I _04073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10361__I0 _04909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07605_ u2.mem\[23\]\[8\] _02913_ _02914_ u2.mem\[22\]\[8\] _03076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08585_ _03811_ u2.mem\[11\]\[5\] _03862_ _03864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06190__B1 _01680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09959__S _04734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07536_ u2.mem\[39\]\[7\] _02855_ _02856_ u2.mem\[48\]\[7\] _03008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08863__S _04033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06447__I _01923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11861__I0 _05903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07467_ u2.mem\[53\]\[6\] _02806_ _02807_ u2.mem\[56\]\[6\] _02940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09206_ _04260_ u2.mem\[25\]\[4\] _04261_ _04262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06418_ _01918_ _01919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07398_ _02868_ _02869_ _02870_ _02871_ _02872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09806__I0 _04570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09137_ _04217_ _00381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06349_ u2.mem\[184\]\[4\] _01778_ _01749_ _01852_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06182__I _01688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09068_ _04176_ _04177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07993__A1 _03441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08019_ _03479_ _03480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_151_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09493__I _04440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11030_ _05386_ u2.mem\[139\]\[2\] _05395_ _05398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08103__S _03546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold1_I output_active_trans.data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11528__I _05667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08793__I0 _03912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12981_ _00860_ clknet_leaf_31_clock u2.mem\[53\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11932_ _05949_ _05960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_3555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10352__I0 _04900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06705__C1 _02092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11863_ _05907_ u2.mem\[191\]\[1\] _05918_ _05920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10814_ _05260_ _01015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08773__S _03978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11794_ _05876_ u2.mem\[186\]\[5\] _05865_ _05877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13533_ _01412_ clknet_leaf_318_clock u2.mem\[192\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10745_ _05218_ u2.mem\[61\]\[10\] _05214_ _05219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10808__S _05253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06484__A1 _01969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07681__B1 _03084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13464_ _01343_ clknet_leaf_344_clock u2.mem\[180\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06484__B2 _01972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10676_ _05175_ _00962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12415_ _00294_ clknet_leaf_160_clock u2.mem\[18\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11604__I0 _05758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07028__A3 _02392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13395_ _01274_ clknet_leaf_307_clock u2.mem\[169\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07188__I _02558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12346_ _00225_ clknet_leaf_59_clock u2.mem\[13\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_179_clock_I clknet_5_30_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06787__A2 _02156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12277_ _00156_ clknet_leaf_102_clock u2.mem\[9\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11907__I1 _03531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11228_ _05523_ _01166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07736__A1 u2.mem\[32\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07736__B2 u2.mem\[2\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11159_ _05478_ _01142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08948__S _04089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13115__CLK clknet_5_22_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_231_clock_I clknet_5_24_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10343__I0 _04891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13265__CLK clknet_leaf_295_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06711__A2 _02126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08370_ _03731_ _00100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07321_ _02470_ _02796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09578__I _04173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06475__A1 _01962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07252_ u2.mem\[18\]\[2\] _02606_ _02608_ u2.mem\[19\]\[2\] _02729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08482__I _03656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07672__B1 _03067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06203_ _01709_ _01710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07183_ _02532_ _02661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07019__A3 _02383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07098__I _02417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06227__A1 u2.mem\[193\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06134_ _01573_ _01574_ _01548_ _01641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_145_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11549__S _05722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06778__A2 _02257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06065_ _01567_ _01571_ _01572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10453__S _05040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08775__I0 _03937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11348__I _05597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09824_ _04596_ u2.mem\[39\]\[9\] _04649_ _04651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06967_ _02432_ _02446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09755_ _04609_ u2.mem\[37\]\[13\] _04606_ _04610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08527__I0 _03829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08706_ _03941_ _03942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08657__I _03663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09686_ _04558_ _00589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10334__I0 _04920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06898_ _02352_ _02376_ _02377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07561__I _02476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08637_ _03824_ u2.mem\[12\]\[11\] _03890_ _03894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11039__A1 _04334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06177__I _01683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08568_ _03831_ u2.mem\[10\]\[14\] _03851_ _03854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12632__CLK clknet_leaf_104_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07519_ _02974_ _02980_ _02985_ _02990_ _02991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_70_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08499_ _03810_ _00150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10530_ _05014_ u2.mem\[56\]\[9\] _05083_ _05085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10262__A2 _04863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10427__I _03717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10461_ _05029_ _05045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_109_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12782__CLK clknet_leaf_253_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12200_ _00079_ clknet_leaf_65_clock u2.mem\[4\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_180_clock_I clknet_5_30_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07415__B1 _02888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13180_ _01059_ clknet_leaf_275_clock u2.mem\[133\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10392_ _04138_ _05000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11762__A2 _05847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12131_ _01472_ clknet_leaf_35_clock u2.driver_mem\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10363__S _04976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13138__CLK clknet_leaf_314_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12062_ data_in_trans\[6\].A clknet_leaf_302_clock data_in_trans\[6\].data_sync vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07718__A1 u2.mem\[26\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08766__I0 _03928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11013_ _05386_ u2.mem\[138\]\[2\] _05382_ _05387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08768__S _03973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07733__A4 _03201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13288__CLK clknet_leaf_364_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12964_ _00843_ clknet_leaf_109_clock u2.mem\[52\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10325__I0 _04911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11915_ _05903_ u2.mem\[193\]\[0\] _05950_ _05951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12895_ _00774_ clknet_leaf_225_clock u2.mem\[48\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09599__S _04506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11846_ _05908_ _01399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11777_ _04287_ _05847_ _05865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11721__I _03666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13516_ _01395_ clknet_leaf_338_clock u2.mem\[189\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10728_ _05004_ _05207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10659_ _05117_ u2.mem\[59\]\[10\] _05162_ _05165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13447_ _01326_ clknet_leaf_343_clock u2.mem\[178\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06209__A1 u2.mem\[152\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10005__A2 _04760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06209__B2 u2.mem\[148\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13378_ _01257_ clknet_leaf_36_clock u2.mem\[166\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12329_ _00208_ clknet_leaf_125_clock u2.mem\[12\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06550__I _02034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07972__A4 _03435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11168__I _05483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07709__B2 u2.mem\[46\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08757__I0 _03919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12505__CLK clknet_leaf_163_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07870_ _03332_ _03333_ _03334_ _03335_ _03336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_110_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10564__I0 _05106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07185__A2 _02515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06821_ u2.mem\[185\]\[4\] _02121_ _02123_ u2.mem\[173\]\[4\] _02302_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06932__A2 _02403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09540_ _04469_ u2.mem\[33\]\[2\] _04465_ _04470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06752_ u2.mem\[146\]\[2\] _02155_ _02157_ u2.mem\[186\]\[2\] _02235_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10316__I0 _04902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07381__I _02618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09182__I0 _04174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12655__CLK clknet_leaf_223_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09471_ _04373_ u2.mem\[31\]\[7\] _04424_ _04428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06683_ u2.mem\[170\]\[1\] _02146_ _02148_ u2.mem\[156\]\[1\] _02167_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08422_ _03689_ u2.mem\[7\]\[7\] _03759_ _03763_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06696__A1 u2.mem\[164\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06696__B2 u2.mem\[178\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08353_ _03718_ _03719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10448__S _05035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09485__I1 u2.mem\[31\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07304_ _01808_ _02361_ _02758_ _02779_ _01495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06448__A1 u2.mem\[193\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11292__I1 u2.mem\[155\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08284_ _03662_ _03663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06448__B2 u2.mem\[194\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09101__I _04181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06999__A2 _02475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07235_ u2.mem\[49\]\[2\] _02660_ _02661_ u2.mem\[46\]\[2\] _02712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12035__CLK clknet_2_3__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07166_ _02640_ _02641_ _02642_ _02643_ _02644_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_117_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11279__S _05545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06117_ u2.mem\[167\]\[0\] _01622_ _01623_ u2.mem\[183\]\[0\] _01624_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07097_ u2.mem\[26\]\[0\] _02573_ _02575_ u2.mem\[10\]\[0\] _02576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07412__A3 _02884_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06048_ _01554_ _01555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12185__CLK clknet_leaf_59_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08748__I0 _03910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13430__CLK clknet_5_4_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09807_ _04641_ _00627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07999_ _01665_ _03462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06923__A2 _02380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10710__I _04986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09738_ _04596_ u2.mem\[37\]\[9\] _04593_ _04597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10307__I0 _04893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_127_clock_I clknet_5_15_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09173__I0 _04161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09669_ _04543_ _04549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11700_ _05817_ _05818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12680_ _00559_ clknet_leaf_129_clock u2.mem\[34\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09212__S _04261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11631_ _05775_ _01317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09476__I1 u2.mem\[31\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06439__A1 u2.mem\[193\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11562_ _05711_ u2.mem\[172\]\[1\] _05731_ _05733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06439__B2 u2.mem\[194\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13301_ _01180_ clknet_leaf_2_clock u2.mem\[153\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10513_ _05075_ _00899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_324_clock clknet_5_7_0_clock clknet_leaf_324_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_13_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11493_ _05689_ _01265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09228__I1 u2.mem\[25\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13232_ _01111_ clknet_leaf_279_clock u2.mem\[142\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10444_ _05001_ u2.mem\[54\]\[4\] _05035_ _05036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08987__I0 _04044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11189__S _05492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13163_ _01042_ clknet_leaf_274_clock u2.mem\[130\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10375_ _04986_ _04987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10794__I0 _05225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12114_ _01477_ clknet_leaf_333_clock u2.select_mem_row\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13094_ _00973_ clknet_leaf_23_clock u2.mem\[60\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11917__S _05950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12024__D mem_address_trans\[9\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12045_ net5 clknet_2_2__leaf_clock_a col_select_trans\[4\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06914__A2 _02391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09164__I0 _04148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07134__C _02394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12947_ _00826_ clknet_leaf_233_clock u2.mem\[51\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08911__I0 _04046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06678__A1 _02049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12878_ _00757_ clknet_leaf_219_clock u2.mem\[47\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10268__S _04923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11829_ _05868_ u2.mem\[189\]\[1\] _05896_ _05898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12058__CLK clknet_leaf_300_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06545__I _02029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_329_clock_I clknet_5_7_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07020_ _02454_ _02496_ _02497_ _02498_ _02499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__06850__A1 u2.mem\[185\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08978__I0 _04035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13453__CLK clknet_leaf_301_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07376__I _02607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10785__I0 _05216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08971_ _04028_ u2.mem\[20\]\[6\] _04102_ _04105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11827__S _05896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07922_ u2.mem\[58\]\[14\] _03275_ _03276_ u2.mem\[36\]\[14\] _03387_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_155_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10537__I0 _05020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07853_ u2.mem\[5\]\[12\] _03153_ _03154_ u2.mem\[38\]\[12\] _03320_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06366__B1 _01721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06905__A2 _02382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06804_ _02277_ _02282_ _02283_ _02284_ _02285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_83_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07784_ _02405_ _03251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09155__I0 _04132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09523_ _04384_ u2.mem\[32\]\[12\] _04458_ _04459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06735_ _02215_ _02216_ _02217_ _02218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11562__S _05731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08902__I0 _04037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09454_ _04417_ _04011_ _04418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06669__A1 u2.mem\[179\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07866__B1 _02448_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06666_ _02150_ _02151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06669__B2 u2.mem\[191\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07330__A2 _02648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08405_ _03480_ _03752_ _03753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_24_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09385_ _04373_ u2.mem\[29\]\[7\] _04367_ _04374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10178__S _04865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06597_ _02081_ _02082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09458__I1 u2.mem\[31\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08336_ _03704_ _03705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08267_ _03572_ u2.mem\[4\]\[12\] _03650_ _03651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09766__I _04617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07218_ u2.mem\[45\]\[2\] _02633_ _02634_ u2.mem\[34\]\[2\] _02695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08670__I _03680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06841__A1 u2.mem\[151\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08198_ _03539_ u2.mem\[3\]\[0\] _03609_ _03610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06841__B2 u2.mem\[158\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08969__I0 _04026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_53_clock_I clknet_5_12_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07149_ _02469_ _02431_ _02433_ _02507_ _02628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_133_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10776__I0 _05207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10160_ _04840_ _04856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_79_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12820__CLK clknet_leaf_61_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11737__S _05840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10091_ _04816_ _00736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10641__S _05152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10528__I0 _05011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12970__CLK clknet_leaf_124_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_278_clock_I clknet_5_21_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12801_ _00680_ clknet_leaf_144_clock u2.mem\[42\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10993_ _05374_ _01080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12732_ _00611_ clknet_leaf_255_clock u2.mem\[38\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13326__CLK clknet_leaf_304_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12663_ _00542_ clknet_leaf_58_clock u2.mem\[33\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_330_clock_I clknet_5_7_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11614_ _05754_ u2.mem\[175\]\[3\] _05761_ _05765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_263_clock clknet_5_23_0_clock clknet_leaf_263_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11256__I1 u2.mem\[153\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12594_ _00473_ clknet_leaf_167_clock u2.mem\[29\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07085__A1 _02451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12019__D net31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12350__CLK clknet_leaf_201_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11545_ _05707_ u2.mem\[171\]\[0\] _05722_ _05723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13476__CLK clknet_leaf_295_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06832__B2 u2.mem\[189\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11476_ _03510_ _05679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13215_ _01094_ clknet_leaf_283_clock u2.mem\[139\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_278_clock clknet_5_21_0_clock clknet_leaf_278_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10427_ _03717_ _05025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10767__I0 _05198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07196__I _02574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10358_ _04977_ _00842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13146_ _01025_ clknet_leaf_38_clock u2.mem\[63\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_5_26_0_clock_I clknet_4_13_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_201_clock clknet_5_28_0_clock clknet_leaf_201_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13077_ _00956_ clknet_leaf_25_clock u2.mem\[59\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10551__S _05095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10289_ _04937_ _00813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10519__I0 _05001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09385__I0 _04373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12028_ row_select_trans\[1\].A clknet_leaf_307_clock row_select_trans\[1\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_7_clock clknet_5_0_0_clock clknet_leaf_7_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_24_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_216_clock clknet_5_28_0_clock clknet_leaf_216_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_81_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06520_ row_select_trans\[5\].data_sync _02005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06451_ _01923_ _01946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07863__A3 _03326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09787__S _04628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09170_ _04237_ _00394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06382_ u2.mem\[167\]\[5\] _01775_ _01776_ u2.mem\[183\]\[5\] _01884_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08121_ _03513_ _03559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07076__A1 _02398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10726__S _05205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08490__I _03667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06823__A1 _02285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08052_ _03507_ _03508_ _03509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12843__CLK clknet_leaf_198_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07003_ _02462_ _02472_ _02478_ _02481_ _02482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_116_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10758__I0 _05227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07379__A2 _02687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08954_ _03629_ _03540_ _03633_ _04094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__12993__CLK clknet_leaf_239_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09376__I0 _04366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07905_ u2.mem\[6\]\[13\] _03327_ _03328_ u2.mem\[47\]\[13\] _03371_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08885_ _04054_ _00292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11183__I0 _05460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07000__A1 _02451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07836_ _02581_ _03303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12223__CLK clknet_leaf_231_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10930__I0 _05305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input16_I data_in_a[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07767_ u2.mem\[23\]\[11\] _03146_ _03147_ u2.mem\[22\]\[11\] _03235_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06894__B _02353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09506_ _04449_ _00518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06718_ u2.mem\[176\]\[1\] _02003_ _02013_ u2.mem\[172\]\[1\] _02019_ u2.mem\[189\]\[1\]
+ _02202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_07698_ u2.mem\[1\]\[10\] _03028_ _03029_ u2.mem\[7\]\[10\] _03167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11486__I1 u2.mem\[167\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07303__A2 _02768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_09437_ _04378_ u2.mem\[30\]\[9\] _04406_ _04408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06649_ _01999_ _02033_ _02134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13499__CLK clknet_leaf_316_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11238__I1 u2.mem\[152\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06185__I _01691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09368_ _04131_ _04362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08319_ data_in_trans\[8\].data_sync _03691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09299_ _04265_ u2.mem\[27\]\[6\] _04318_ _04321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11330_ _05583_ u2.mem\[158\]\[0\] _05585_ _05586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06814__A1 u2.mem\[169\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08106__S _03546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06814__B2 u2.mem\[147\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11261_ _05542_ _01180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10212_ _04885_ u2.mem\[49\]\[0\] _04887_ _04888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13000_ _00879_ clknet_leaf_322_clock u2.mem\[54\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11192_ _05497_ _01156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10143_ _04792_ u2.mem\[47\]\[4\] _04846_ _04847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07790__A2 _03250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10074_ _04804_ u2.mem\[45\]\[9\] _04802_ _04805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11266__I _05545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06750__B1 _02147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12716__CLK clknet_leaf_254_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_10976_ _04224_ _05363_ _05364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_71_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12715_ _00594_ clknet_leaf_252_clock u2.mem\[37\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11930__S _05955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11229__I1 u2.mem\[151\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06095__I _01601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12646_ _00525_ clknet_leaf_93_clock u2.mem\[32\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12866__CLK clknet_leaf_151_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12577_ _00456_ clknet_leaf_170_clock u2.mem\[28\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06805__B2 u2.mem\[189\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11528_ _05667_ _05711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08007__B1 _03462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11459_ _05666_ _01254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_140_clock clknet_5_13_0_clock clknet_leaf_140_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07230__A1 u2.mem\[53\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13129_ _01008_ clknet_leaf_327_clock u2.mem\[62\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07230__B2 u2.mem\[56\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09358__I0 _04285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07654__I _02527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12246__CLK clknet_leaf_73_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input8_I data_in_a[10] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08670_ _03680_ _03917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_155_clock clknet_5_27_0_clock clknet_leaf_155_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_27_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10912__I0 _05301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07621_ _02613_ _03092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12396__CLK clknet_leaf_180_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07552_ u2.mem\[27\]\[8\] _03021_ _03022_ u2.mem\[35\]\[8\] _03023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06503_ row_select_trans\[2\].data_sync _01988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07483_ u2.mem\[9\]\[6\] _02836_ _02837_ u2.mem\[25\]\[6\] _02956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06219__B _01725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09222_ _04272_ u2.mem\[25\]\[9\] _04270_ _04273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06434_ _01923_ _01933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09153_ _04128_ u2.mem\[24\]\[1\] _04226_ _04228_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06365_ u2.mem\[144\]\[4\] _01670_ _01672_ u2.mem\[182\]\[4\] _01868_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_226_clock_I clknet_5_25_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08104_ _03547_ _00018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06257__C1 _01705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09084_ _04140_ u2.mem\[22\]\[4\] _04187_ _04188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11640__I1 u2.mem\[177\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06296_ u2.mem\[170\]\[2\] _01687_ _01689_ u2.mem\[156\]\[2\] _01801_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08035_ _01545_ _03490_ _03495_ _00001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13021__CLK clknet_leaf_258_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09597__I0 _04476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_108_clock clknet_5_11_0_clock clknet_leaf_108_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_107_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07221__A1 u2.mem\[27\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06024__A2 _01517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09986_ _04739_ _04750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_104_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09349__I0 _04276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07772__A2 _03153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13171__CLK clknet_leaf_264_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08937_ _04032_ u2.mem\[19\]\[8\] _04084_ _04085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11156__I0 _05464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08596__S _03867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08868_ _04043_ _00286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10903__I0 _05307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07524__A2 _02993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07819_ _03257_ _03269_ _03278_ _03285_ _03286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_85_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08799_ _03997_ _00263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10830_ _05269_ _01022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10761_ _05229_ u2.mem\[61\]\[15\] _05223_ _05230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11750__S _05849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12500_ _00379_ clknet_leaf_105_clock u2.mem\[23\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13480_ _01359_ clknet_leaf_289_clock u2.mem\[183\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10692_ _05173_ _05184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_8_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12431_ _00310_ clknet_leaf_160_clock u2.mem\[19\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12119__CLK clknet_leaf_332_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12362_ _00241_ clknet_leaf_134_clock u2.mem\[14\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11313_ _05411_ _05566_ _05575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_12293_ _00172_ clknet_leaf_101_clock u2.mem\[10\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12269__CLK clknet_leaf_185_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09588__I0 _04467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11244_ _05511_ u2.mem\[152\]\[3\] _05529_ _05533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06799__B _01993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08260__I0 _03566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11175_ _05468_ u2.mem\[148\]\[3\] _05484_ _05488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07763__A2 _03066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10126_ _04813_ u2.mem\[46\]\[13\] _04835_ _04837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_72_clock clknet_5_8_0_clock clknet_leaf_72_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_95_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11147__I0 _05470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12032__D row_select_trans\[3\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10057_ _04783_ _04793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_114_1565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07515__A2 _02890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_175_clock_I clknet_5_27_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_87_clock clknet_5_11_0_clock clknet_leaf_87_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10370__I1 u2.mem\[52\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11724__I _03670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07142__C _02364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10959_ _05353_ _01067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_10_clock clknet_5_1_0_clock clknet_leaf_10_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_31_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09130__S _04213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06981__C _02364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12629_ _00508_ clknet_leaf_97_clock u2.mem\[31\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13044__CLK clknet_leaf_26_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06150_ _01656_ _01657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_25_clock clknet_5_2_0_clock clknet_leaf_25_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06081_ _01587_ _01588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07451__B2 u2.mem\[47\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09579__I0 _04496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13194__CLK clknet_leaf_272_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09840_ _04224_ _04659_ _04660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08251__I0 _03557_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07384__I _02613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07754__A2 _03049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09771_ _04573_ u2.mem\[38\]\[2\] _04618_ _04621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_06983_ u2.mem\[15\]\[0\] _02457_ _02461_ u2.mem\[13\]\[0\] _02462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11138__I0 _05464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11835__S _05895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08722_ _03921_ u2.mem\[14\]\[7\] _03947_ _03951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11689__I1 u2.mem\[180\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09751__I0 _04605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08653_ _03480_ _03904_ _03905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_113_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07604_ _03065_ _03068_ _03071_ _03074_ _03075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_1609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08584_ _03863_ _00182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06190__A1 u2.mem\[147\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06190__B2 u2.mem\[169\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07535_ u2.mem\[5\]\[7\] _02920_ _02921_ u2.mem\[38\]\[7\] _03007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11570__S _05730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07466_ u2.mem\[54\]\[6\] _02881_ _02882_ u2.mem\[55\]\[6\] _02939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11861__I1 u2.mem\[191\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09040__S _04155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09205_ _04251_ _04261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06417_ _01911_ _01916_ _01918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07690__A1 _03138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07397_ u2.mem\[27\]\[5\] _02788_ _02789_ u2.mem\[35\]\[5\] _02871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09975__S _04740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09136_ _04164_ u2.mem\[23\]\[11\] _04213_ _04217_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06348_ u2.mem\[171\]\[4\] _01611_ _01770_ u2.mem\[157\]\[4\] _01851_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13537__CLK clknet_leaf_14_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09067_ data_in_trans\[15\].data_sync _04176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06279_ _01781_ _01782_ _01783_ _01784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_11_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10914__S _05319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07993__A2 _03446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08018_ _03477_ mem_address_trans\[5\].data_sync _03478_ mem_address_trans\[7\].data_sync
+ _03479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_162_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12561__CLK clknet_leaf_170_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08242__I0 _03548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_8_0_clock clknet_3_4_0_clock clknet_4_8_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_49_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09969_ _04681_ u2.mem\[43\]\[0\] _04740_ _04741_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12980_ _00859_ clknet_leaf_43_clock u2.mem\[53\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09215__S _04261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09742__I0 _04599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11931_ _05959_ _01433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06705__C2 u2.mem\[177\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06638__I _02122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06181__A1 _01566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11862_ _05919_ _01404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09014__I _04134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06720__A3 _02194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10813_ u2.mem\[63\]\[5\] _03511_ _05258_ _05260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13067__CLK clknet_leaf_248_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11301__I0 _05544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11793_ _03679_ _05876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09949__I _04718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13532_ _01411_ clknet_leaf_334_clock u2.mem\[192\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08853__I _04014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10744_ _03700_ _05218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07130__B1 _02608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13463_ _01342_ clknet_leaf_344_clock u2.mem\[180\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06484__A2 _01970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10675_ _05093_ u2.mem\[60\]\[0\] _05174_ _05175_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12414_ _00293_ clknet_leaf_178_clock u2.mem\[18\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12091__CLK clknet_2_3__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13394_ _01273_ clknet_leaf_310_clock u2.mem\[169\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12345_ _00224_ clknet_leaf_60_clock u2.mem\[13\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12027__D net38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10824__S _05263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12276_ _00155_ clknet_leaf_102_clock u2.mem\[9\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11227_ _05508_ u2.mem\[151\]\[2\] _05520_ _05523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07197__B1 _02674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10040__I0 _04716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11158_ _05466_ u2.mem\[147\]\[2\] _05475_ _05478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10109_ _04827_ _00743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11089_ _05434_ _05435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_62_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11454__I _03491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08964__S _04097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06172__A1 _01678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09110__A1 _03752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09859__I _04660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07320_ _02464_ _02795_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12434__CLK clknet_leaf_124_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07251_ u2.mem\[52\]\[2\] _02601_ _02603_ u2.mem\[21\]\[2\] _02728_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07672__A1 u2.mem\[29\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06475__A2 _01955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06202_ _01600_ _01634_ _01709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07182_ _02530_ _02660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06133_ _01639_ _01640_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07424__A1 _02872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12584__CLK clknet_leaf_115_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09594__I _04500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06064_ _01547_ _01570_ _01571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08204__S _03609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11359__I0 _05595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10031__I0 _04707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09823_ _04650_ _00634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09754_ _04608_ _04609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06966_ _02430_ _02445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_86_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08527__I1 u2.mem\[9\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08705_ _03607_ _03726_ _03878_ _03941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_67_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09685_ _04489_ u2.mem\[36\]\[11\] _04554_ _04558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11364__I _05607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06897_ _02341_ _02342_ _02376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08636_ _03893_ _00204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06163__A1 _01638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08567_ _03853_ _00175_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07518_ _02986_ _02987_ _02988_ _02989_ _02990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08673__I _03684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08498_ _03808_ u2.mem\[9\]\[4\] _03809_ _03810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07449_ u2.mem\[39\]\[5\] _02855_ _02856_ u2.mem\[48\]\[5\] _02923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_126_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10460_ _05044_ _00877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11598__I0 _05754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_123_clock_I clknet_5_15_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09119_ _04207_ _00373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06218__A2 _01669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10391_ _04999_ _00853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_159_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10270__I0 _04893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12130_ _01471_ clknet_leaf_35_clock u2.driver_mem\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07966__A2 _03427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10443__I _05029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12061_ net19 clknet_2_0__leaf_clock_a data_in_trans\[6\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07718__A2 _03139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09009__I _04130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10022__I0 _04698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09963__I0 _04714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11012_ _05342_ _05386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12307__CLK clknet_leaf_104_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11770__I0 _05833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12963_ _00842_ clknet_leaf_109_clock u2.mem\[52\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11914_ _05949_ _05950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_73_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12457__CLK clknet_leaf_126_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12894_ _00773_ clknet_leaf_214_clock u2.mem\[48\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_48_clock_I clknet_5_7_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11845_ _05907_ u2.mem\[190\]\[1\] _05905_ _05908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11776_ _03655_ _05864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13515_ _01394_ clknet_leaf_340_clock u2.mem\[189\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10727_ _05206_ _00982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13446_ _01325_ clknet_leaf_350_clock u2.mem\[177\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10658_ _05164_ _00955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11589__I0 _05746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10554__S _05095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13377_ _01256_ clknet_leaf_11_clock u2.mem\[166\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10589_ _03713_ _05124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12328_ _00207_ clknet_leaf_126_clock u2.mem\[12\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10961__A1 _05354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12259_ _00138_ clknet_leaf_70_clock u2.mem\[8\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10013__I0 _04689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07709__A2 _03126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09954__I0 _04705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11385__S _05616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_325_clock_I clknet_5_7_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13232__CLK clknet_leaf_279_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06820_ u2.mem\[144\]\[4\] _02115_ _02117_ u2.mem\[182\]\[4\] _02301_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06393__A1 u2.mem\[166\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06393__B2 u2.mem\[161\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07662__I _02558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06932__A3 _02392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06751_ u2.mem\[179\]\[2\] _02150_ _02152_ u2.mem\[191\]\[2\] _02234_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11513__I0 _05668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09470_ _04427_ _00504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06682_ u2.mem\[185\]\[1\] _02121_ _02123_ u2.mem\[173\]\[1\] _02166_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08694__S _03933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08421_ _03762_ _00120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10729__S _05205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07893__B2 u2.mem\[11\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08493__I _03671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08352_ _03717_ _03718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07303_ _02763_ _02768_ _02773_ _02778_ _02779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__06448__A2 _01942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08283_ _03496_ _03662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07234_ u2.mem\[14\]\[2\] _02657_ _02658_ u2.mem\[12\]\[2\] _02711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07165_ u2.mem\[3\]\[1\] _02480_ _02359_ _02643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_145_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10464__S _05045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06116_ _01571_ _01617_ _01623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06605__C1 u2.mem\[193\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08070__A1 _03521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07096_ _02574_ _02575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_160_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10263__I _04922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06047_ _01553_ _01554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06620__A2 _02104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09945__I0 _04696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11752__I0 _05829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09806_ _04570_ u2.mem\[39\]\[1\] _04639_ _04641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06384__A1 u2.mem\[184\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07572__I _02499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07998_ _01547_ _03461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09737_ _04595_ _04596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06949_ _02427_ _02428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09668_ _04548_ _00581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08619_ _03806_ u2.mem\[12\]\[3\] _03880_ _03884_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10639__S _05152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09599_ _04478_ u2.mem\[34\]\[6\] _04506_ _04509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07884__B2 u2.mem\[20\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11630_ _05754_ u2.mem\[176\]\[3\] _05771_ _05775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08109__S _03546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08684__I0 _03926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11561_ _05732_ _01290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13300_ _01179_ clknet_leaf_2_clock u2.mem\[153\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10512_ _04992_ u2.mem\[56\]\[1\] _05073_ _05075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13105__CLK clknet_leaf_314_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11492_ _05680_ u2.mem\[167\]\[5\] _05682_ _05689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_274_clock_I clknet_5_21_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13231_ _01110_ clknet_leaf_284_clock u2.mem\[142\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08436__I0 _03715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10443_ _05029_ _05035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_136_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08987__I1 u2.mem\[20\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13162_ _01041_ clknet_leaf_275_clock u2.mem\[130\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10374_ _04117_ _04986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11269__I _05504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10794__I1 u2.mem\[62\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10173__I _04864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12113_ _01476_ clknet_leaf_331_clock u2.select_mem_row\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13255__CLK clknet_leaf_295_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13093_ _00972_ clknet_leaf_24_clock u2.mem\[60\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09936__I0 _04687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12044_ col_select_trans\[3\].A clknet_leaf_299_clock col_select_trans\[3\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11743__I0 _05835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_5_0_clock clknet_0_clock clknet_3_5_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_133_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06914__A3 _02392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09164__I1 u2.mem\[24\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12946_ _00825_ clknet_leaf_233_clock u2.mem\[51\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06127__A1 _01549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06678__A2 _02074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12877_ _00756_ clknet_leaf_214_clock u2.mem\[47\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11828_ _05897_ _01392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11997__CLK clknet_leaf_33_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07627__A1 _03064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11759_ _05854_ _01366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08427__I0 _03698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10284__S _04933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13429_ _01308_ clknet_leaf_337_clock u2.mem\[175\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06850__A2 _02120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07657__I _02532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10234__I0 _04902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08978__I1 u2.mem\[20\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08052__A1 _03507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11982__I0 _05225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10083__I _04783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08970_ _04104_ _00327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07921_ u2.mem\[53\]\[14\] _03272_ _03273_ u2.mem\[56\]\[14\] _03386_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12622__CLK clknet_leaf_189_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07852_ _03309_ _03312_ _03315_ _03318_ _03319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_84_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07392__I _02443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06366__B2 u2.mem\[185\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06905__A3 _02383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06803_ u2.mem\[165\]\[4\] _02076_ _02079_ u2.mem\[163\]\[4\] u2.mem\[145\]\[4\]
+ _02082_ _02284_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_56_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput1 col_select_a[0] net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07783_ u2.mem\[32\]\[12\] _03248_ _03249_ u2.mem\[2\]\[12\] _03250_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09522_ _04442_ _04458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12772__CLK clknet_leaf_91_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06734_ u2.mem\[159\]\[2\] _02174_ _02176_ u2.mem\[149\]\[2\] _02217_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06118__A1 _01586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09453_ _04416_ _04417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_149_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06665_ _01998_ _02077_ _02150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10459__S _05040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_08404_ _03751_ _03752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_5_7_0_clock clknet_4_3_0_clock clknet_5_7_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_101_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09384_ _04150_ _04373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12002__CLK clknet_leaf_42_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06596_ _02044_ _02080_ _02081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_5_0_0_clock_I clknet_4_0_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08335_ data_in_trans\[11\].data_sync _03704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08266_ _03634_ _03650_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07217_ _01726_ _02361_ _02665_ _02694_ _01493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12152__CLK clknet_leaf_64_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08418__I0 _03681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10194__S _04875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13278__CLK clknet_leaf_9_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08197_ _03608_ _03609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_106_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10225__I0 _04895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08969__I1 u2.mem\[20\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08043__A1 _01769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07148_ _02626_ _02627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11089__I _05434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10776__I1 u2.mem\[62\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11973__I0 _05216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07079_ _02551_ _02537_ _02538_ _02442_ _02558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__10922__S _05327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10090_ _04815_ u2.mem\[45\]\[14\] _04811_ _04816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11725__I0 _05833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07149__A3 _02433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10721__I _04997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12800_ _00679_ clknet_leaf_144_clock u2.mem\[42\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07306__B1 _02634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10992_ _05335_ u2.mem\[137\]\[0\] _05373_ _05374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_76_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12731_ _00610_ clknet_leaf_216_clock u2.mem\[38\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12662_ _00541_ clknet_leaf_76_clock u2.mem\[33\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06646__I _02130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11613_ _05764_ _01310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12593_ _00472_ clknet_leaf_167_clock u2.mem\[29\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10464__I0 _05023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07085__A2 _02452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11544_ _05721_ _05722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_51_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06293__B1 _01701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08409__I0 _03664_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11475_ _05678_ _01258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13214_ _01093_ clknet_leaf_282_clock u2.mem\[139\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08034__A1 _03492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10426_ _05024_ _00863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11964__I0 _05915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11928__S _05955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12035__D net42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13145_ _01024_ clknet_leaf_39_clock u2.mem\[63\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10357_ _04904_ u2.mem\[52\]\[8\] _04976_ _04977_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06596__A1 _02044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09909__I0 _04703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08302__S _03677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13076_ _00955_ clknet_leaf_24_clock u2.mem\[59\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10288_ _04911_ u2.mem\[50\]\[11\] _04933_ _04937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11716__I0 _05825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11727__I _03674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12795__CLK clknet_leaf_220_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12027_ net38 clknet_2_0__leaf_clock_a row_select_trans\[1\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06348__A1 u2.mem\[171\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06348__B2 u2.mem\[157\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12025__CLK clknet_2_3__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07848__A1 u2.mem\[52\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12929_ _00808_ clknet_leaf_233_clock u2.mem\[50\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06450_ u2.mem\[0\]\[6\] _01945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_107_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12175__CLK clknet_leaf_218_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06381_ u2.mem\[178\]\[5\] _01772_ _01773_ u2.mem\[164\]\[5\] _01883_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13420__CLK clknet_leaf_298_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08120_ _03558_ _00023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10455__I0 _05014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08051_ _03493_ _03508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06823__A2 _02290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07387__I _02623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10207__I0 _04817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07002_ u2.mem\[3\]\[0\] _02480_ _02359_ _02481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13570__CLK clknet_leaf_14_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11955__I0 _05907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08820__I0 _03939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10742__S _05214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08953_ _04093_ _00321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11707__I0 _05794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11637__I _05778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07904_ u2.mem\[8\]\[13\] _03324_ _03325_ u2.mem\[4\]\[13\] _03370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08884_ _04019_ u2.mem\[18\]\[2\] _04051_ _04054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06339__A1 _01809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11183__I1 u2.mem\[149\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_222_clock_I clknet_5_28_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07835_ _02579_ _03302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07000__A2 _02452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_323_clock clknet_5_18_0_clock clknet_leaf_323_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07766_ _03230_ _03231_ _03232_ _03233_ _03234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_37_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07850__I _02607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09505_ _04366_ u2.mem\[32\]\[4\] _04448_ _04449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06717_ u2.mem\[194\]\[1\] _02198_ _02199_ u2.mem\[190\]\[1\] _02200_ u2.mem\[160\]\[1\]
+ _02201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_38_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12518__CLK clknet_leaf_94_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07697_ u2.mem\[15\]\[10\] _03025_ _03026_ u2.mem\[13\]\[10\] _03166_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07303__A3 _02773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_09436_ _04407_ _00490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08882__S _04051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06648_ _01992_ _02052_ _02133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_338_clock clknet_5_5_0_clock clknet_leaf_338_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_52_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_09367_ _04361_ _00467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06579_ _02057_ _02064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10446__I0 _05005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08318_ _03690_ _00089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09298_ _04320_ _00439_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12668__CLK clknet_leaf_193_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08249_ _03554_ u2.mem\[4\]\[4\] _03640_ _03641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06814__A2 _02142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11260_ _05514_ u2.mem\[153\]\[4\] _05536_ _05542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11946__I0 _05227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10211_ _04886_ _04887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10652__S _05157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08811__I0 _03930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11191_ _05470_ u2.mem\[149\]\[4\] _05491_ _05497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06578__A1 u2.mem\[167\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07775__B1 _03095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06578__B2 u2.mem\[183\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10142_ _04840_ _04846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08122__S _03555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10073_ _04595_ _04804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08856__I _03697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06750__A1 u2.mem\[170\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06750__B2 u2.mem\[156\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10099__S _04820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12198__CLK clknet_leaf_73_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10975_ _05275_ _05363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__13443__CLK clknet_leaf_356_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_12714_ _00593_ clknet_leaf_49_clock u2.mem\[36\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06376__I _01877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12645_ _00524_ clknet_leaf_93_clock u2.mem\[32\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09687__I _04543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10437__I0 _04992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08591__I _03856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12576_ _00455_ clknet_leaf_169_clock u2.mem\[28\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10626__I _05130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11527_ _05710_ _01278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_171_clock_I clknet_5_27_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11458_ _05663_ u2.mem\[166\]\[0\] _05665_ _05666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11937__I0 _05218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10409_ _05011_ u2.mem\[53\]\[8\] _05012_ _05013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08802__I0 _03921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06569__A1 _02052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11389_ _05595_ u2.mem\[161\]\[5\] _05615_ _05622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13128_ _01007_ clknet_leaf_46_clock u2.mem\[62\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07230__A2 _02486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13059_ _00938_ clknet_leaf_27_clock u2.mem\[58\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06995__B _02384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07620_ _02611_ _03091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07670__I _02574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06741__A1 u2.mem\[144\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06741__B2 u2.mem\[182\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_31_0_clock clknet_4_15_0_clock clknet_5_31_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07551_ _02435_ _03022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_96_clock_I clknet_5_10_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09798__S _04633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06502_ _01985_ _01986_ _01987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07482_ u2.mem\[29\]\[6\] _02833_ _02834_ u2.mem\[11\]\[6\] _02955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09221_ _04157_ _04272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12810__CLK clknet_leaf_139_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06433_ u2.mem\[192\]\[2\] _01931_ _01932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10428__I0 _05025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09152_ _04227_ _00386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06364_ u2.mem\[154\]\[4\] _01699_ _01701_ u2.mem\[162\]\[4\] _01866_ _01867_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_147_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08207__S _03614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08103_ _03539_ u2.mem\[1\]\[0\] _03546_ _03547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06257__C2 u2.mem\[194\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09083_ _04181_ _04187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06295_ u2.mem\[173\]\[2\] _01720_ _01722_ u2.mem\[185\]\[2\] _01800_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10536__I _05072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08034_ _03492_ _03494_ _03495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11928__I0 _05209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11568__S _05730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09597__I1 u2.mem\[34\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10472__S _05051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07757__B1 _03133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10600__I0 _05093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07221__A2 _02428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13316__CLK clknet_leaf_300_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09985_ _04749_ _00697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08936_ _04073_ _04084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_135_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11156__I1 u2.mem\[147\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_262_clock clknet_5_23_0_clock clknet_leaf_262_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_135_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08867_ _04041_ u2.mem\[17\]\[12\] _04042_ _04043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12340__CLK clknet_leaf_80_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13466__CLK clknet_leaf_347_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07818_ _03279_ _03280_ _03281_ _03284_ _03285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_17_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08676__I _03688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08798_ _03917_ u2.mem\[16\]\[5\] _03995_ _03997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06732__A1 u2.mem\[187\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06732__B2 u2.mem\[192\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07749_ u2.mem\[58\]\[11\] _03042_ _03043_ u2.mem\[36\]\[11\] _03217_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_277_clock clknet_5_21_0_clock clknet_leaf_277_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06196__I _01702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07288__A2 _02673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10760_ _03721_ _05229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12490__CLK clknet_leaf_121_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09419_ _04360_ u2.mem\[30\]\[1\] _04396_ _04398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_4_4_0_clock clknet_3_2_0_clock clknet_4_4_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_10691_ _05183_ _00969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_200_clock clknet_5_28_0_clock clknet_leaf_200_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12430_ _00309_ clknet_leaf_178_clock u2.mem\[19\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06924__I _02402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11092__I0 _05424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12361_ _00240_ clknet_leaf_133_clock u2.mem\[14\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06799__A1 u2.mem\[184\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11312_ _05574_ _01199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12292_ _00171_ clknet_leaf_101_clock u2.mem\[10\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_215_clock clknet_5_28_0_clock clknet_leaf_215_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_153_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11919__I0 _05909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11243_ _05532_ _01172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10382__S _04989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07748__B1 _03040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07212__A2 _02617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11174_ _05487_ _01148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08260__I1 u2.mem\[4\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10125_ _04836_ _00750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08787__S _03990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11147__I1 u2.mem\[146\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10056_ _04578_ _04792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06723__A1 u2.mem\[167\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_118_clock_I clknet_5_15_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06723__B2 u2.mem\[183\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07920__B1 _02511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12833__CLK clknet_leaf_148_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07279__A2 _02660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10958_ _05352_ u2.mem\[134\]\[5\] _05336_ _05353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10557__S _05095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10889_ _05307_ u2.mem\[130\]\[5\] _05296_ _05308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12983__CLK clknet_leaf_326_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12628_ _00507_ clknet_leaf_97_clock u2.mem\[31\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09276__I0 _04281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10356__I _04965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11083__I0 _05430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12559_ _00438_ clknet_leaf_170_clock u2.mem\[27\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12213__CLK clknet_leaf_68_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06080_ _01550_ _01579_ _01587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_89_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13339__CLK clknet_leaf_4_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08400__A1 _03605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08251__I1 u2.mem\[4\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09770_ _04620_ _00611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08697__S _03933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06982_ _02460_ _02461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_1543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08721_ _03950_ _00232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08496__I _03675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10897__I0 _05301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08652_ _03903_ _03904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_94_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07603_ u2.mem\[28\]\[8\] _03072_ _03073_ u2.mem\[31\]\[8\] _03074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08583_ _03808_ u2.mem\[11\]\[4\] _03862_ _03863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06190__A2 _01676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11851__S _05905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07534_ _03002_ _03003_ _03004_ _03005_ _03006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_78_1494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06478__B1 _01948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07465_ u2.mem\[50\]\[6\] _02878_ _02879_ u2.mem\[51\]\[6\] _02938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09204_ _04139_ _04260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06416_ _01916_ _01917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09267__I0 _04272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07396_ u2.mem\[40\]\[5\] _02785_ _02786_ u2.mem\[30\]\[5\] _02870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07690__A2 _03145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09120__I _04202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09135_ _04216_ _00380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09967__A1 _04311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11074__I0 _05424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06347_ u2.mem\[167\]\[4\] _01775_ _01776_ u2.mem\[183\]\[4\] _01850_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07978__B1 _02575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09066_ _04175_ _00352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06278_ u2.mem\[172\]\[2\] _01654_ _01667_ u2.mem\[150\]\[2\] _01783_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06650__B1 _02134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08017_ mem_address_trans\[6\].data_sync _03478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07993__A3 _03451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12706__CLK clknet_leaf_238_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09991__S _04750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08242__I1 u2.mem\[4\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06402__B1 _01688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09968_ _04739_ _04740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10930__S _05326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08919_ _04010_ u2.mem\[19\]\[0\] _04074_ _04075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12856__CLK clknet_leaf_129_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09899_ _04696_ u2.mem\[41\]\[6\] _04692_ _04697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11930_ _05211_ u2.mem\[193\]\[7\] _05955_ _05959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06919__I _02363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06705__A1 u2.mem\[165\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07902__B1 _02629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06705__B2 u2.mem\[163\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11861_ _05903_ u2.mem\[191\]\[0\] _05918_ _05919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06181__A2 _01629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10812_ _05259_ _01014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06720__A4 _02203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11792_ _05875_ _01378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11301__I1 u2.mem\[156\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06469__B1 _01943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13531_ _01410_ clknet_leaf_333_clock u2.mem\[192\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10743_ _05217_ _00987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12236__CLK clknet_leaf_211_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13462_ _01341_ clknet_leaf_346_clock u2.mem\[180\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09258__I0 _04263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07681__A2 _03083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10674_ _05173_ _05174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09030__I _04147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12413_ _00292_ clknet_leaf_197_clock u2.mem\[18\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13393_ _01272_ clknet_5_16_0_clock u2.mem\[169\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_154_clock clknet_5_27_0_clock clknet_leaf_154_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07969__B1 _02533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12344_ _00223_ clknet_leaf_131_clock u2.mem\[13\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12386__CLK clknet_leaf_224_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_44_clock_I clknet_5_6_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12275_ _00154_ clknet_leaf_102_clock u2.mem\[9\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11226_ _05522_ _01165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09430__I0 _04371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_169_clock clknet_5_27_0_clock clknet_leaf_169_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07197__A1 u2.mem\[26\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12043__D net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11157_ _05477_ _01141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06944__A1 _02422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10108_ _04795_ u2.mem\[46\]\[5\] _04825_ _04827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11088_ _04417_ _05402_ _05434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_48_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10039_ _04780_ _00720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_269_clock_I clknet_5_22_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09205__I _04251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13011__CLK clknet_leaf_323_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_107_clock clknet_5_11_0_clock clknet_leaf_107_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_63_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09141__S _04218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07121__A1 _02547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07250_ u2.mem\[17\]\[2\] _02591_ _02593_ u2.mem\[24\]\[2\] _02727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09249__I0 _04254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08980__S _04107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_321_clock_I clknet_5_18_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07672__A2 _03066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13161__CLK clknet_leaf_276_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11056__I0 _05380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06201_ _01707_ _01708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07181_ u2.mem\[14\]\[1\] _02657_ _02658_ u2.mem\[12\]\[1\] _02659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12729__CLK clknet_leaf_44_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06132_ _01638_ _01576_ _01639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07424__A2 _02877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06063_ _01569_ _01570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11359__I1 u2.mem\[159\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12879__CLK clknet_leaf_230_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09421__I0 _04362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09822_ _04592_ u2.mem\[39\]\[8\] _04649_ _04650_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06935__A1 _02407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09753_ data_in_trans\[13\].data_sync _04608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06965_ _02443_ _02444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08220__S _03619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12109__CLK clknet_leaf_140_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08704_ _03940_ _00225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09684_ _04557_ _00588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06148__C1 u2.mem\[172\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06896_ _02374_ _02375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_67_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08635_ _03822_ u2.mem\[12\]\[10\] _03890_ _03893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06163__A2 _01634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08566_ _03829_ u2.mem\[10\]\[13\] _03851_ _03853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12259__CLK clknet_leaf_70_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13504__CLK clknet_leaf_331_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07517_ u2.mem\[43\]\[7\] _02816_ _02817_ u2.mem\[20\]\[7\] _02989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08497_ _03799_ _03809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_35_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08160__I0 _03548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07448_ u2.mem\[5\]\[5\] _02920_ _02921_ u2.mem\[38\]\[5\] _02922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_71_clock clknet_5_8_0_clock clknet_leaf_71_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_11_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11047__I0 _05388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07379_ u2.mem\[5\]\[4\] _02687_ _02688_ u2.mem\[38\]\[4\] _02854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_13_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11598__I1 u2.mem\[174\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09118_ _04136_ u2.mem\[23\]\[3\] _04203_ _04207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07415__A2 _02887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06218__A3 _01724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10390_ _04998_ u2.mem\[53\]\[3\] _04989_ _04999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09049_ _04162_ _00348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_86_clock clknet_5_11_0_clock clknet_leaf_86_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_89_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10724__I _05000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12060_ data_in_trans\[5\].A clknet_leaf_300_clock data_in_trans\[5\].data_sync vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11756__S _05849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11011_ _05385_ _01087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06926__A1 _02398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06387__C1 _01577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11770__I1 u2.mem\[185\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13034__CLK clknet_leaf_326_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12962_ _00841_ clknet_leaf_156_clock u2.mem\[52\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_270_clock_I clknet_5_20_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09025__I _04143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11913_ _04013_ _05926_ _05949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_4099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_24_clock clknet_5_2_0_clock clknet_leaf_24_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12893_ _00772_ clknet_leaf_214_clock u2.mem\[48\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11844_ _03662_ _05907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11286__I0 _05544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11775_ _05863_ _01373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08151__I0 _03579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11986__A1 _03535_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13514_ _01393_ clknet_leaf_340_clock u2.mem\[189\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10726_ _05204_ u2.mem\[61\]\[4\] _05205_ _05206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_39_clock clknet_5_6_0_clock clknet_leaf_39_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_144_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_1_0_clock clknet_0_clock clknet_3_1_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_158_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13445_ _01324_ clknet_leaf_350_clock u2.mem\[177\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10657_ _05115_ u2.mem\[59\]\[9\] _05162_ _05164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11589__I1 u2.mem\[174\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13376_ _01255_ clknet_leaf_10_clock u2.mem\[166\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10588_ _05123_ _00926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12327_ _00206_ clknet_leaf_126_clock u2.mem\[12\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06090__A1 _01576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12258_ _00137_ clknet_leaf_228_clock u2.mem\[8\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11209_ _03502_ _05510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12189_ _00068_ clknet_leaf_252_clock u2.mem\[4\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09136__S _04213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06393__A2 _01592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06750_ u2.mem\[170\]\[2\] _02145_ _02147_ u2.mem\[156\]\[2\] _02233_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06559__I _02022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12401__CLK clknet_leaf_161_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13527__CLK clknet_leaf_316_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06681_ u2.mem\[144\]\[1\] _02115_ _02117_ u2.mem\[182\]\[1\] _02165_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08420_ _03685_ u2.mem\[7\]\[6\] _03759_ _03762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_0_0_clock_I clknet_3_0_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08351_ data_in_trans\[14\].data_sync _03717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12551__CLK clknet_leaf_115_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08142__I0 _03572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07302_ _02774_ _02775_ _02776_ _02777_ _02778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06508__B _01992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08282_ _03661_ _00082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07233_ u2.mem\[44\]\[2\] _02654_ _02655_ u2.mem\[42\]\[2\] _02710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06853__B1 _02157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10745__S _05214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07164_ u2.mem\[16\]\[1\] _02475_ _02477_ u2.mem\[33\]\[1\] _02642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06115_ _01571_ _01607_ _01622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_173_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06605__C2 _02089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07095_ _02566_ _02567_ _02493_ _02568_ _02574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__08070__A2 _03519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06046_ _01547_ _01549_ _01552_ _01553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_5_3_0_clock clknet_4_1_0_clock clknet_5_3_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_114_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11576__S _05739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13057__CLK clknet_leaf_240_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09945__I1 u2.mem\[42\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06908__A1 _02365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11752__I1 u2.mem\[184\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09805_ _04640_ _00626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input39_I row_select_a[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07997_ u2.active_mem\[4\] _03458_ _03459_ u2.active_mem\[5\] _03460_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_101_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06948_ _02418_ _02420_ _02425_ _02426_ _02427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_09736_ data_in_trans\[9\].data_sync _04595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09667_ _04471_ u2.mem\[36\]\[3\] _04544_ _04548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06879_ _02357_ _02358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08618_ _03883_ _00196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09598_ _04508_ _00551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08549_ _03843_ _00167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07097__B1 _02575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11560_ _05707_ u2.mem\[172\]\[0\] _05731_ _05732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10511_ _05074_ _00898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06844__B1 _02116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10655__S _05162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11491_ _05688_ _01264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_217_clock_I clknet_5_28_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13230_ _01109_ clknet_leaf_279_clock u2.mem\[141\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10442_ _05034_ _00869_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08125__S _03555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13161_ _01040_ clknet_leaf_276_clock u2.mem\[130\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10373_ _04985_ _00849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12112_ _01475_ clknet_leaf_334_clock u2.select_mem_row\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13092_ _00971_ clknet_leaf_24_clock u2.mem\[60\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11486__S _05683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12043_ net4 clknet_2_2__leaf_clock_a col_select_trans\[3\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10390__S _04989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08859__I _03701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11743__I1 u2.mem\[183\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12424__CLK clknet_leaf_123_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11285__I _05558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12945_ _00824_ clknet_leaf_233_clock u2.mem\[51\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07875__A2 _03338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12876_ _00755_ clknet_leaf_215_clock u2.mem\[47\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06678__A3 _02113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11827_ _05864_ u2.mem\[189\]\[0\] _05896_ _05897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07627__A2 _03075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11758_ _05835_ u2.mem\[184\]\[4\] _05848_ _05854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08824__A1 _03483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10709_ _05193_ _00977_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11689_ _05790_ u2.mem\[180\]\[1\] _05810_ _05812_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13428_ _01307_ clknet_leaf_350_clock u2.mem\[174\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_2_0__f_clock_a clknet_0_clock_a clknet_2_0__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_31_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13359_ _01238_ clknet_leaf_357_clock u2.mem\[163\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07260__B1 _02715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07920_ u2.mem\[54\]\[14\] _02509_ _02511_ u2.mem\[55\]\[14\] _03385_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07851_ u2.mem\[18\]\[12\] _03316_ _03317_ u2.mem\[19\]\[12\] _03318_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11195__I _03491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06366__A2 _01719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06802_ u2.mem\[188\]\[4\] _02185_ _02186_ u2.mem\[187\]\[4\] _02187_ u2.mem\[192\]\[4\]
+ _02283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__12917__CLK clknet_leaf_83_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07782_ _02395_ _03249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput2 col_select_a[1] net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09521_ _04457_ _00525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06733_ u2.mem\[188\]\[2\] _02185_ _02177_ u2.mem\[175\]\[2\] _02216_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07315__A1 u2.mem\[27\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06118__A2 _01617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11923__I _05949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_166_clock_I clknet_5_26_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09452_ _03748_ _03902_ _04416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06664_ u2.mem\[170\]\[0\] _02146_ _02148_ u2.mem\[156\]\[0\] _02149_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07866__A2 _02444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_08403_ _03748_ _03750_ _03751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09383_ _04372_ _00472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06595_ _01991_ _02017_ _02080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08334_ _03703_ _00092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08265_ _03649_ _00077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_4_0_clock_I clknet_4_2_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07216_ _02672_ _02679_ _02686_ _02693_ _02694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_165_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09615__I0 _04494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08196_ _03605_ _03606_ _03483_ _03607_ _03608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_146_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07147_ _02458_ _02459_ _02484_ _02364_ _02626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_161_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_26_0_clock clknet_4_13_0_clock clknet_5_26_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_145_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11973__I1 u2.mem\[194\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07251__B1 _02603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12447__CLK clknet_leaf_159_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07078_ u2.mem\[57\]\[0\] _02554_ _02556_ u2.mem\[41\]\[0\] _02557_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_126_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06029_ u2.driver_mem\[12\] _01517_ _01537_ _01520_ _01538_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_133_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08679__I _03692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11725__I1 u2.mem\[182\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07149__A4 _02507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09719_ _04143_ _04582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10991_ _05372_ _05373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_74_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07306__A1 u2.mem\[45\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08354__I0 _03719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12730_ _00609_ clknet_leaf_43_clock u2.mem\[37\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06927__I _02405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10161__I0 _04810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09303__I _04312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12661_ _00540_ clknet_leaf_77_clock u2.mem\[33\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08106__I0 _03548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11612_ _05752_ u2.mem\[175\]\[2\] _05761_ _05764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12592_ _00471_ clknet_leaf_168_clock u2.mem\[29\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11543_ _04310_ _05690_ _05721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_106_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13222__CLK clknet_leaf_280_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06293__A1 u2.mem\[154\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09606__I0 _04485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06293__B2 u2.mem\[162\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11474_ _05677_ u2.mem\[166\]\[4\] _05664_ _05678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13213_ _01092_ clknet_leaf_282_clock u2.mem\[139\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11413__I0 _05623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10425_ _05023_ u2.mem\[53\]\[13\] _05021_ _05024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11964__I1 u2.mem\[194\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07242__B1 _02556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13144_ _01023_ clknet_leaf_39_clock u2.mem\[63\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10356_ _04965_ _04976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__13372__CLK clknet_leaf_359_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06596__A2 _02080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13075_ _00954_ clknet_leaf_25_clock u2.mem\[59\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10287_ _04936_ _00812_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11716__I1 u2.mem\[182\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12026_ row_select_trans\[0\].A clknet_leaf_302_clock row_select_trans\[0\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06330__C _01833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11944__S _05965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12051__D net14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10152__I0 _04801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12928_ _00807_ clknet_leaf_235_clock u2.mem\[50\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12859_ _00738_ clknet_leaf_199_clock u2.mem\[46\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06380_ _01879_ _01880_ _01881_ _01882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10295__S _04938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08050_ _03506_ _03507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07481__B1 _02907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06572__I _02006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06284__B2 u2.mem\[161\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06823__A3 _02303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07001_ _02479_ _02480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06036__A1 u3.data vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07233__B1 _02655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11955__I1 u2.mem\[194\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_92_clock_I clknet_5_10_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08952_ _04048_ u2.mem\[19\]\[15\] _04089_ _04093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11707__I1 u2.mem\[181\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07903_ u2.mem\[39\]\[13\] _03321_ _03322_ u2.mem\[48\]\[13\] _03369_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08883_ _04053_ _00291_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11854__S _05904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07834_ u2.mem\[29\]\[12\] _03299_ _03300_ u2.mem\[11\]\[12\] _03301_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07765_ u2.mem\[28\]\[11\] _03072_ _03073_ u2.mem\[31\]\[11\] _03233_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09504_ _04442_ _04448_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06716_ _02137_ _02200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07696_ _03161_ _03162_ _03163_ _03164_ _03165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10143__I0 _04792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09435_ _04375_ u2.mem\[30\]\[8\] _04406_ _04407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06647_ u2.mem\[148\]\[0\] _02129_ _02131_ u2.mem\[152\]\[0\] _02132_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13245__CLK clknet_leaf_285_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_09366_ _04360_ u2.mem\[29\]\[1\] _04358_ _04361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06578_ u2.mem\[167\]\[0\] _02060_ _02062_ u2.mem\[183\]\[0\] _02063_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_1556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08317_ _03689_ u2.mem\[5\]\[7\] _03677_ _03690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09297_ _04263_ u2.mem\[27\]\[5\] _04318_ _04320_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07578__I _02514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07472__B1 _02894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08248_ _03634_ _03640_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_126_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13395__CLK clknet_leaf_307_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08179_ _03597_ _00043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09793__I _04617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10210_ _04013_ _04863_ _04886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07224__B1 _02471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11190_ _05496_ _01155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10141_ _04845_ _00757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_0_0_clock clknet_3_0_0_clock clknet_4_0_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_10072_ _04803_ _00730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11764__S _05857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10382__I0 _04992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06750__A2 _02145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06657__I _02141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10134__I0 _04782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10974_ _05362_ _01073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09033__I data_in_trans\[7\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_56_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12713_ _00592_ clknet_leaf_50_clock u2.mem\[36\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09968__I _04739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12644_ _00523_ clknet_leaf_92_clock u2.mem\[32\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08872__I _03718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11634__I0 _05758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12575_ _00454_ clknet_leaf_183_clock u2.mem\[28\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10907__I _05318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06266__A1 u2.mem\[171\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06266__B2 u2.mem\[157\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11526_ _05707_ u2.mem\[170\]\[0\] _05709_ _05710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_114_clock_I clknet_5_14_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12046__D col_select_trans\[4\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08007__A2 _03461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11457_ _05664_ _05665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10843__S _05278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12762__CLK clknet_5_13_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11937__I1 u2.mem\[193\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10408_ _04988_ _05012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_67_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11388_ _05621_ _01228_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06569__A2 _02053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10339_ _04885_ u2.mem\[52\]\[0\] _04966_ _04967_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13127_ _01006_ clknet_leaf_327_clock u2.mem\[62\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09208__I _04144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13058_ _00937_ clknet_leaf_242_clock u2.mem\[58\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08566__I0 _03829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11674__S _05801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12009_ net26 clknet_2_0__leaf_clock_a mem_address_trans\[2\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06995__C _02473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12142__CLK clknet_leaf_211_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11473__I _05676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13268__CLK clknet_leaf_9_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07550_ _02427_ _03021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_39_clock_I clknet_5_6_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06501_ row_select_trans\[1\].data_sync _01986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07481_ u2.mem\[26\]\[6\] _02906_ _02907_ u2.mem\[10\]\[6\] _02954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07297__A3 _02771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09220_ _04271_ _00410_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06432_ _01919_ _01931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08782__I mem_address_trans\[7\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12292__CLK clknet_leaf_101_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09151_ _04119_ u2.mem\[24\]\[0\] _04226_ _04227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06363_ _01863_ _01864_ _01865_ _01866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10428__I1 u2.mem\[53\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08102_ _03545_ _03546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_148_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06257__A1 u2.mem\[190\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09082_ _04186_ _00357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07454__B1 _02898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11250__A1 _04248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06294_ u2.mem\[144\]\[2\] _01671_ _01673_ u2.mem\[182\]\[2\] _01799_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08033_ _03493_ _03494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07206__B1 _02603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09984_ _04698_ u2.mem\[43\]\[7\] _04745_ _04749_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08935_ _04083_ _00313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08557__I0 _03820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11584__S _05738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_316_clock_I clknet_5_18_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08957__I _04096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08866_ _04014_ _04042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_3706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07861__I _02623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input21_I data_in_a[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07817_ u2.mem\[43\]\[12\] _03282_ _03283_ u2.mem\[20\]\[12\] _03284_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_3739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08797_ _03996_ _00262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_5_12_0_clock_I clknet_4_6_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09989__S _04750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11069__A1 _04394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07748_ u2.mem\[53\]\[11\] _03039_ _03040_ u2.mem\[56\]\[11\] _03216_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07679_ u2.mem\[17\]\[9\] _03077_ _03078_ u2.mem\[24\]\[9\] _03149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10928__S _05327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06496__A1 _01981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09418_ _04397_ _00482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08692__I _03709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10690_ _05110_ u2.mem\[60\]\[7\] _05179_ _05183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11616__I0 _05756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09349_ _04276_ u2.mem\[28\]\[11\] _04346_ _04350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12785__CLK clknet_leaf_235_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12360_ _00239_ clknet_leaf_136_clock u2.mem\[14\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07101__I _02579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11311_ _05556_ u2.mem\[156\]\[5\] _05567_ _05574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12291_ _00170_ clknet_leaf_103_clock u2.mem\[10\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12015__CLK clknet_2_2__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11919__I1 u2.mem\[193\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11242_ _05508_ u2.mem\[152\]\[2\] _05529_ _05532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06940__I _02389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08796__I0 _03914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11173_ _05466_ u2.mem\[148\]\[2\] _05484_ _05487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10124_ _04810_ u2.mem\[46\]\[12\] _04835_ _04836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06420__A1 u2.mem\[193\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06420__B2 u2.mem\[192\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12165__CLK clknet_leaf_91_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08548__I0 _03811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10055_ _04791_ _00725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13410__CLK clknet_leaf_305_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_40_clock_I clknet_5_6_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13560__CLK clknet_leaf_32_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10957_ _05351_ _05352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08720__I0 _03919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11480__A1 _05354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10888_ _05004_ _05307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12627_ _00506_ clknet_leaf_97_clock u2.mem\[31\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12558_ _00437_ clknet_leaf_191_clock u2.mem\[27\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07987__A1 _03447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_265_clock_I clknet_5_23_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_322_clock clknet_5_18_0_clock clknet_leaf_322_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_145_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11509_ _04248_ _05690_ _05699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_12489_ _00368_ clknet_leaf_121_clock u2.mem\[22\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09139__S _04218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08787__I0 _03900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11468__I _03502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12508__CLK clknet_leaf_180_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08978__S _04107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_337_clock clknet_5_4_0_clock clknet_leaf_337_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_101_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_06981_ _02458_ _02459_ _02442_ _02364_ _02460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08539__I0 _03802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13090__CLK clknet_leaf_242_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08720_ _03919_ u2.mem\[14\]\[6\] _03947_ _03950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11299__A1 _04333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12658__CLK clknet_leaf_224_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08651_ _03901_ _03902_ _03903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07602_ _02586_ _03073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07911__B2 u2.mem\[30\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08582_ _03856_ _03862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_26_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07533_ u2.mem\[18\]\[7\] _02850_ _02851_ u2.mem\[19\]\[7\] _03005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_78_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10748__S _05214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08711__I0 _03910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06478__A1 u2.mem\[193\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07464_ _02933_ _02934_ _02935_ _02936_ _02937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08218__S _03619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09401__I _04357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09203_ _04259_ _00405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06415_ _01912_ _01916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10547__I _05094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07395_ u2.mem\[32\]\[5\] _02782_ _02783_ u2.mem\[2\]\[5\] _02869_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09267__I1 u2.mem\[26\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07690__A3 _03152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09134_ _04161_ u2.mem\[23\]\[10\] _04213_ _04216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12038__CLK clknet_leaf_302_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06346_ u2.mem\[178\]\[4\] _01772_ _01773_ u2.mem\[164\]\[4\] _01849_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07427__B1 _02900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09967__A2 _04659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08017__I mem_address_trans\[6\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07978__B2 u2.mem\[10\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09065_ _04174_ u2.mem\[21\]\[14\] _04168_ _04175_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06277_ u2.mem\[174\]\[2\] _01657_ _01658_ u2.mem\[155\]\[2\] _01661_ u2.mem\[181\]\[2\]
+ _01782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__10483__S _05056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08016_ mem_address_trans\[4\].data_sync _03477_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06650__A1 u2.mem\[194\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06650__B2 u2.mem\[190\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07993__A4 _03456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12188__CLK clknet_leaf_252_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11378__I _05615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13433__CLK clknet_leaf_338_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09967_ _04311_ _04659_ _04739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_103_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08918_ _04073_ _04074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_135_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09898_ _04585_ _04696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07591__I _02555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08849_ _03688_ _04030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08950__I0 _04046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11860_ _05917_ _05918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11837__I0 _05876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10811_ u2.mem\[63\]\[4\] _03507_ _05258_ _05259_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11791_ _05874_ u2.mem\[186\]\[4\] _05865_ _05875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11841__I _05904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06469__A1 u2.mem\[193\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13530_ _01409_ clknet_leaf_317_clock u2.mem\[191\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06469__B2 u2.mem\[194\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10742_ _05216_ u2.mem\[61\]\[9\] _05214_ _05217_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07130__A2 _02606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13461_ _01340_ clknet_leaf_344_clock u2.mem\[180\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10673_ _04334_ _05172_ _05173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09258__I1 u2.mem\[26\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12412_ _00291_ clknet_leaf_198_clock u2.mem\[18\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07418__B1 _02891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13392_ _01271_ clknet_leaf_353_clock u2.mem\[168\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12343_ _00222_ clknet_leaf_132_clock u2.mem\[13\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12274_ _00153_ clknet_leaf_166_clock u2.mem\[9\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11225_ _05505_ u2.mem\[151\]\[1\] _05520_ _05522_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08798__S _03995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07197__A2 _02673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11156_ _05464_ u2.mem\[147\]\[1\] _05475_ _05477_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06944__A2 _02350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10107_ _04826_ _00742_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10328__I0 _04913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11087_ _05433_ _01115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10038_ _04714_ u2.mem\[44\]\[14\] _04777_ _04780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08941__I0 _04037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12950__CLK clknet_leaf_30_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06172__A3 _01588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_0_0_clock_I clknet_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11989_ _00001_ clknet_leaf_318_clock u2.mem\[0\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09221__I _04157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13306__CLK clknet_leaf_358_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07121__A2 _02371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09249__I1 u2.mem\[26\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06200_ _01556_ _01677_ _01593_ _01707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__07409__B1 _02882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07180_ _02527_ _02658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_261_clock clknet_5_23_0_clock clknet_leaf_261_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_118_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06131_ _01557_ _01638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_157_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12330__CLK clknet_leaf_125_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13456__CLK clknet_leaf_304_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07424__A3 _02886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07676__I _02595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06062_ _01558_ _01568_ _01569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11198__I _05501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_276_clock clknet_5_21_0_clock clknet_leaf_276_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_160_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09421__I1 u2.mem\[30\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10567__I0 _05108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12480__CLK clknet_leaf_164_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09821_ _04638_ _04649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_113_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06396__B1 _01709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06935__A2 _02408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09752_ _04607_ _00606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06964_ _02398_ _02438_ _02439_ _02442_ _02443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__10319__I0 _04904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08703_ _03939_ u2.mem\[13\]\[15\] _03933_ _03940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08300__I _03675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06895_ _02373_ _02374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09683_ _04487_ u2.mem\[36\]\[10\] _04554_ _04557_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06148__C2 _01654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08932__I0 _04028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08634_ _03892_ _00203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_5_clock clknet_5_0_0_clock clknet_leaf_5_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_214_clock clknet_5_28_0_clock clknet_leaf_214_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_82_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11819__I0 _05872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08565_ _03852_ _00174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10478__S _05051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07516_ u2.mem\[49\]\[7\] _02893_ _02894_ u2.mem\[46\]\[7\] _02988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08496_ _03675_ _03808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08160__I1 u2.mem\[2\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07447_ _02628_ _02921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06320__B1 _01635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_229_clock clknet_5_25_0_clock clknet_leaf_229_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_13_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06871__A1 col_select_trans\[5\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07378_ _02843_ _02846_ _02849_ _02852_ _02853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_104_1533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09117_ _04206_ _00372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06329_ _01830_ _01831_ _01832_ _01833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_8_clock_I clknet_5_1_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09048_ _04161_ u2.mem\[21\]\[10\] _04155_ _04162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07820__B1 _03133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12823__CLK clknet_leaf_135_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11010_ _05384_ u2.mem\[138\]\[1\] _05382_ _05385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06387__C2 u2.mem\[193\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_1545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_213_clock_I clknet_5_29_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12961_ _00840_ clknet_leaf_157_clock u2.mem\[52\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08923__I0 _04019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11912_ _01981_ _05929_ _05948_ _01425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07887__B1 _02561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12892_ _00771_ clknet_leaf_209_clock u2.mem\[48\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12203__CLK clknet_leaf_217_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13329__CLK clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11843_ _05906_ _01398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07270__B _02745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11286__I1 u2.mem\[155\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11774_ _05837_ u2.mem\[185\]\[5\] _05856_ _05863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13513_ _01392_ clknet_leaf_340_clock u2.mem\[189\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11986__A2 _05972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10725_ _05195_ _05205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12353__CLK clknet_leaf_150_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13479__CLK clknet_leaf_290_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06862__A1 col_select_trans\[5\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13444_ _01323_ clknet_leaf_349_clock u2.mem\[177\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10656_ _05163_ _00954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10587_ _05121_ u2.mem\[57\]\[12\] _05122_ _05123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13375_ _01254_ clknet_leaf_352_clock u2.mem\[166\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12326_ _00205_ clknet_leaf_85_clock u2.mem\[12\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12054__D data_in_trans\[2\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06090__A2 _01596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12257_ _00136_ clknet_leaf_228_clock u2.mem\[8\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10851__S _05277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09417__S _04396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11208_ _05509_ _01160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12188_ _00067_ clknet_leaf_252_clock u2.mem\[4\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06378__C2 u2.mem\[181\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11139_ _05465_ _01135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11682__S _05800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06680_ u2.mem\[169\]\[1\] _02142_ _02144_ u2.mem\[147\]\[1\] _02164_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11481__I _05682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08350_ _03716_ _00095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11426__A1 _04094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07301_ u2.mem\[6\]\[3\] _02622_ _02624_ u2.mem\[47\]\[3\] _02777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08281_ _03657_ u2.mem\[5\]\[0\] _03660_ _03661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07232_ _02705_ _02706_ _02707_ _02708_ _02709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_clkbuf_4_4_0_clock_I clknet_3_2_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06853__A1 u2.mem\[146\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06853__B2 u2.mem\[186\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12846__CLK clknet_leaf_203_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07163_ u2.mem\[1\]\[1\] _02465_ _02471_ u2.mem\[7\]\[1\] _02641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06605__A1 u2.mem\[151\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06114_ u2.mem\[178\]\[0\] _01618_ _01620_ u2.mem\[164\]\[0\] _01621_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07094_ _02572_ _02573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_162_clock_I clknet_5_26_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06605__B2 u2.mem\[158\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11857__S _05904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06045_ _01550_ _01551_ _01552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12996__CLK clknet_leaf_33_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09327__S _04336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06369__B1 _01693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09804_ _04565_ u2.mem\[39\]\[0\] _04639_ _04640_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10560__I _05094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12226__CLK clknet_leaf_143_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07996_ _01613_ _03459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09735_ _04594_ _00602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06947_ _02412_ _02426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11592__S _05748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_153_clock clknet_5_25_0_clock clknet_leaf_153_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_28_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09666_ _04547_ _00580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06878_ _02347_ _02351_ _02356_ _02357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_82_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08617_ _03804_ u2.mem\[12\]\[2\] _03880_ _03883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_5_22_0_clock clknet_4_11_0_clock clknet_5_22_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09597_ _04476_ u2.mem\[34\]\[5\] _04506_ _04508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11391__I _05499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_87_clock_I clknet_5_11_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07090__B _02425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08548_ _03811_ u2.mem\[10\]\[5\] _03841_ _03843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_168_clock clknet_5_27_0_clock clknet_leaf_168_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_23_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08479_ _03796_ _00144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06844__A1 u2.mem\[144\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10510_ _04987_ u2.mem\[56\]\[0\] _05073_ _05074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11490_ _05677_ u2.mem\[167\]\[4\] _05682_ _05688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06844__B2 u2.mem\[182\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10441_ _04998_ u2.mem\[54\]\[3\] _05030_ _05034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10372_ _04920_ u2.mem\[52\]\[15\] _04981_ _04985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13160_ _01039_ clknet_leaf_276_clock u2.mem\[130\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07939__A4 _03403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12111_ _01474_ clknet_leaf_332_clock u2.select_mem_row\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13001__CLK clknet_leaf_322_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13091_ _00970_ clknet_leaf_22_clock u2.mem\[60\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12042_ col_select_trans\[2\].A clknet_leaf_299_clock col_select_trans\[2\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_106_clock clknet_5_11_0_clock clknet_leaf_106_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_105_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_364_clock_I clknet_5_0_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12719__CLK clknet_leaf_236_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08875__I _03722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12944_ _00823_ clknet_leaf_235_clock u2.mem\[51\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12875_ _00754_ clknet_leaf_218_clock u2.mem\[47\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06678__A4 _02162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11007__S _05382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11826_ _05895_ _05896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12869__CLK clknet_leaf_80_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09700__S _04567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12049__D net7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11757_ _05853_ _01365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07627__A3 _03086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06835__A1 u2.mem\[187\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10708_ _05128_ u2.mem\[60\]\[15\] _05189_ _05193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06835__B2 u2.mem\[192\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11688_ _05811_ _01338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13427_ _01306_ clknet_leaf_349_clock u2.mem\[174\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10645__I _05151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10639_ _05097_ u2.mem\[59\]\[1\] _05152_ _05154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08115__I _03545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13358_ _01237_ clknet_leaf_356_clock u2.mem\[163\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12309_ _00188_ clknet_leaf_100_clock u2.mem\[11\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07260__A1 _01768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13289_ _01168_ clknet_leaf_1_clock u2.mem\[151\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12249__CLK clknet_leaf_55_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11476__I _03510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10380__I _04126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07850_ _02607_ _03317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10942__I0 _05340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_70_clock clknet_5_8_0_clock clknet_leaf_70_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06801_ u2.mem\[171\]\[4\] _02066_ _02068_ u2.mem\[157\]\[4\] _02281_ _02282_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_116_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07781_ _02385_ _03248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12399__CLK clknet_leaf_155_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06771__B1 _02067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput3 col_select_a[2] net3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09520_ _04382_ u2.mem\[32\]\[11\] _04453_ _04457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06732_ u2.mem\[187\]\[2\] _02186_ _02187_ u2.mem\[192\]\[2\] _02215_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_109_clock_I clknet_5_11_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09560__I0 _04482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09451_ _04415_ _00497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06663_ _02147_ _02148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_85_clock clknet_5_11_0_clock clknet_leaf_85_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_36_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08402_ _03749_ _03632_ _03750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09382_ _04371_ u2.mem\[29\]\[6\] _04367_ _04372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06594_ _02078_ _02079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09610__S _04511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07079__A1 _02551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08333_ _03702_ u2.mem\[5\]\[10\] _03694_ _03703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08264_ _03570_ u2.mem\[4\]\[11\] _03645_ _03649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06826__A1 u2.mem\[164\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07215_ _02689_ _02690_ _02691_ _02692_ _02693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08195_ _03541_ _03607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_140_1563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07146_ u2.mem\[6\]\[0\] _02622_ _02624_ u2.mem\[47\]\[0\] _02625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_5_8_0_clock_I clknet_4_4_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_23_clock clknet_5_2_0_clock clknet_leaf_23_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_156_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07077_ _02555_ _02556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09379__I0 _04369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13174__CLK clknet_leaf_275_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06028_ u2.driver_mem\[13\] _01518_ _01537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_121_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10290__I _04922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07085__B _02442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_38_clock clknet_5_6_0_clock clknet_leaf_38_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_101_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07979_ u2.mem\[29\]\[15\] _03299_ _03300_ u2.mem\[11\]\[15\] _03443_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_19_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09718_ _04581_ _00598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10990_ _04249_ _05363_ _05372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_55_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07306__A2 _02633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09649_ _04521_ _04537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_16_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12660_ _00539_ clknet_leaf_75_clock u2.mem\[33\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09520__S _04453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11611_ _05763_ _01309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12591_ _00470_ clknet_leaf_172_clock u2.mem\[29\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11110__I0 _05426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06817__A1 u2.mem\[148\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11542_ _05720_ _01283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07490__A1 _02959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06293__A2 _01699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11473_ _05676_ _05677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13212_ _01091_ clknet_leaf_291_clock u2.mem\[138\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10424_ _03713_ _05023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11413__I1 u2.mem\[163\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13517__CLK clknet_leaf_318_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11497__S _05692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13143_ _01022_ clknet_leaf_39_clock u2.mem\[63\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10355_ _04975_ _00841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07242__B2 u2.mem\[41\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10286_ _04909_ u2.mem\[50\]\[10\] _04933_ _04936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13074_ _00953_ clknet_leaf_241_clock u2.mem\[59\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11177__I0 _05470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12541__CLK clknet_leaf_188_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12025_ net37 clknet_2_3__leaf_clock_a row_select_trans\[0\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10924__I0 _05299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08742__A1 _03605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_110_clock_I clknet_5_14_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12927_ _00806_ clknet_leaf_234_clock u2.mem\[50\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11960__S _05975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06339__B _01842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12858_ _00737_ clknet_leaf_129_clock u2.mem\[45\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11809_ _05885_ _01385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13047__CLK clknet_leaf_44_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12789_ _00668_ clknet_leaf_71_clock u2.mem\[41\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06808__A1 u2.mem\[155\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06808__B2 u2.mem\[150\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07076__A4 _02552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10375__I _04986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07481__B2 u2.mem\[10\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07000_ _02451_ _02452_ _02434_ _02455_ _02479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__12071__CLK clknet_2_1__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_35_clock_I clknet_5_3_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08281__I0 _03657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08951_ _04092_ _00320_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07902_ u2.mem\[5\]\[13\] _02627_ _02629_ u2.mem\[38\]\[13\] _03368_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08882_ _04017_ u2.mem\[18\]\[1\] _04051_ _04053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07833_ _02569_ _03300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07764_ u2.mem\[9\]\[11\] _03069_ _03070_ u2.mem\[25\]\[11\] _03232_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09404__I _04170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09503_ _04447_ _00517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06715_ _02134_ _02199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07695_ u2.mem\[27\]\[10\] _03021_ _03022_ u2.mem\[35\]\[10\] _03164_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09434_ _04395_ _04406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_53_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06646_ _02130_ _02131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09365_ _04127_ _04360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06577_ _02061_ _02062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08316_ _03688_ _03689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_312_clock_I clknet_5_17_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09296_ _04319_ _00438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08247_ _03639_ _00069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08178_ _03566_ u2.mem\[2\]\[9\] _03595_ _03597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07129_ _02607_ _02608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11110__S _05445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07775__A2 _03094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10140_ _04790_ u2.mem\[47\]\[3\] _04841_ _04845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06983__B1 _02461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10071_ _04801_ u2.mem\[45\]\[8\] _04802_ _04803_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11859__A1 _04416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11844__I _03662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10382__I1 u2.mem\[53\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06938__I _02387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10973_ _05352_ u2.mem\[135\]\[5\] _05355_ _05362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12712_ _00591_ clknet_leaf_50_clock u2.mem\[36\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07160__B1 _02436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12643_ _00522_ clknet_leaf_94_clock u2.mem\[32\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12094__CLK clknet_leaf_218_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06673__I _02157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12574_ _00453_ clknet_leaf_186_clock u2.mem\[28\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10598__A1 _04288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11525_ _05708_ _05709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_141_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12907__CLK clknet_leaf_221_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11456_ _04179_ _05645_ _05664_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_32_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10407_ _03691_ _05011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11387_ _05593_ u2.mem\[161\]\[4\] _05615_ _05621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13126_ _01005_ clknet_leaf_23_clock u2.mem\[62\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10338_ _04965_ _04966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_112_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11955__S _05972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12062__D data_in_trans\[6\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13057_ _00936_ clknet_leaf_240_clock u2.mem\[58\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10269_ _04926_ _00804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08566__I1 u2.mem\[10\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09763__I0 _04615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12008_ mem_address_trans\[1\].A clknet_leaf_299_clock mem_address_trans\[1\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11570__I0 _05719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_261_clock_I clknet_5_23_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09224__I _04160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06500_ _01984_ _01985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07480_ _02949_ _02950_ _02951_ _02952_ _02953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07151__B1 _02629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06431_ _01727_ _01915_ _01926_ _01930_ _01465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09150_ _04225_ _04226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_148_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06583__I _02067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06362_ u2.mem\[152\]\[4\] _01713_ _01715_ u2.mem\[148\]\[4\] _01865_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08101_ _03483_ _03542_ _03544_ _03545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_30_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07454__A1 _01877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09081_ _04136_ u2.mem\[22\]\[3\] _04182_ _04186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06293_ u2.mem\[154\]\[2\] _01699_ _01701_ u2.mem\[162\]\[2\] _01797_ _01798_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_163_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08032_ _03488_ _03493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11389__I0 _05595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10061__I0 _04795_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07757__A2 _03132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09983_ _04748_ _00696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08934_ _04030_ u2.mem\[19\]\[7\] _04079_ _04083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08865_ _03709_ _04041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11664__I _05676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13212__CLK clknet_leaf_291_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07816_ _02516_ _03283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08796_ _03914_ u2.mem\[16\]\[4\] _03995_ _03996_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06193__A1 _01615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input14_I data_in_a[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07747_ u2.mem\[54\]\[11\] _03114_ _03115_ u2.mem\[55\]\[11\] _03215_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07678_ u2.mem\[23\]\[9\] _03146_ _03147_ u2.mem\[22\]\[9\] _03148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_13_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13362__CLK clknet_leaf_354_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_5_16_0_clock_I clknet_4_8_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09417_ _04356_ u2.mem\[30\]\[0\] _04396_ _04397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07693__A1 u2.mem\[32\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06629_ _02045_ _02002_ _02114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06496__A2 _01927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09348_ _04349_ _00460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11616__I1 u2.mem\[175\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07445__A1 _02915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09279_ _04308_ _00432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11310_ _05573_ _01198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12290_ _00169_ clknet_leaf_165_clock u2.mem\[10\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11839__I _03655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11241_ _05531_ _01171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07748__A2 _03039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09993__I0 _04707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11172_ _05486_ _01147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10123_ _04819_ _04835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_121_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06420__A2 _01917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08548__I1 u2.mem\[10\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10054_ _04790_ u2.mem\[45\]\[3\] _04784_ _04791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06668__I _02152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06184__A1 _01566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07920__A2 _02509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10956_ _04143_ _05351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08720__I1 u2.mem\[14\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06487__A2 _01917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11480__A2 _05645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10887_ _05306_ _01042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12626_ _00505_ clknet_leaf_170_clock u2.mem\[31\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07436__A1 u2.mem\[9\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12057__D net17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07436__B2 u2.mem\[25\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12557_ _00436_ clknet_leaf_192_clock u2.mem\[27\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_208_clock_I clknet_5_29_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10291__I0 _04913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11508_ _05698_ _01271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12488_ _00367_ clknet_leaf_164_clock u2.mem\[22\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11749__I _05848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11439_ _05653_ _01247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09984__I0 _04698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11791__I0 _05874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13235__CLK clknet_leaf_272_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13109_ _00988_ clknet_leaf_19_clock u2.mem\[61\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06980_ _02419_ _02459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_101_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09155__S _04226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input6_I col_select_a[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09361__A1 _03904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08650_ _03749_ _03877_ _03902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07601_ _02584_ _03072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13385__CLK clknet_leaf_306_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08581_ _03861_ _00181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07532_ u2.mem\[52\]\[7\] _02847_ _02848_ u2.mem\[21\]\[7\] _03004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07463_ u2.mem\[3\]\[6\] _02801_ _02745_ _02936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06478__A2 _01960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10828__I _05252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09202_ _04258_ u2.mem\[25\]\[3\] _04252_ _04259_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06414_ _01914_ _01915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07394_ u2.mem\[45\]\[5\] _02866_ _02867_ u2.mem\[34\]\[5\] _02868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07202__I _02595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07690__A4 _03159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09133_ _04215_ _00379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07427__A1 u2.mem\[61\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06345_ _01845_ _01846_ _01847_ _01848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07978__A2 _02573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10282__I0 _04904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09064_ _04173_ _04174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06276_ u2.mem\[189\]\[2\] _01649_ _01663_ u2.mem\[180\]\[2\] _01651_ u2.mem\[176\]\[2\]
+ _01781_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_162_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08015_ u3.data _03476_ net43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08227__I0 _03575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06650__A2 _02133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10563__I _05004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09129__I _04202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10034__I0 _04709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09975__I0 _04689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08033__I _03493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11595__S _05748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11782__I0 _05868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06402__A2 _01686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09966_ _04738_ _00689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12602__CLK clknet_leaf_113_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08917_ _04072_ _03988_ _04073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_4205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09897_ _04695_ _00663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07093__B _02493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08848_ _04029_ _00280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07902__A2 _02627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_4_clock_I clknet_5_0_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08779_ _03486_ _03983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_166_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_157_clock_I clknet_5_26_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12752__CLK clknet_leaf_227_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10810_ _05252_ _05258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07115__B1 _02593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11837__I1 u2.mem\[189\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11790_ _03674_ _05874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06469__A2 _01960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10738__I _05195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10741_ _03696_ _05216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13460_ _01339_ clknet_leaf_345_clock u2.mem\[180\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10672_ _04862_ _05172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13108__CLK clknet_leaf_20_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07112__I _02590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12411_ _00290_ clknet_leaf_177_clock u2.mem\[18\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07418__B2 u2.mem\[12\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13391_ _01270_ clknet_leaf_353_clock u2.mem\[168\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07969__A2 _02531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10273__I0 _04895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12342_ _00221_ clknet_leaf_78_clock u2.mem\[13\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08091__A1 _01980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08218__I0 _03566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13258__CLK clknet_leaf_312_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12132__CLK clknet_leaf_34_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12273_ _00152_ clknet_leaf_165_clock u2.mem\[9\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06641__A2 _02125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09039__I _04123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10025__I0 _04700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_5_17_0_clock clknet_4_8_0_clock clknet_5_17_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_11224_ _05521_ _01164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11155_ _05476_ _01140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07782__I _02395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12282__CLK clknet_leaf_119_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10106_ _04792_ u2.mem\[46\]\[4\] _04825_ _04826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11086_ _05432_ u2.mem\[142\]\[5\] _05421_ _05433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10037_ _04779_ _00719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10849__S _05278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11988_ _00000_ clknet_leaf_362_clock u3.data vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10939_ _05338_ _01062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_4_0_clock_I clknet_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08118__I _03511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_12609_ _00488_ clknet_leaf_155_clock u2.mem\[30\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_359_clock_I clknet_5_1_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10264__I0 _04885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06130_ u2.mem\[188\]\[0\] _01631_ _01633_ u2.mem\[187\]\[0\] _01636_ u2.mem\[192\]\[0\]
+ _01637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_173_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08082__A1 _01969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07424__A4 _02897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08209__I0 _03557_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06061_ col_select_trans\[3\].data_sync _01568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10016__I0 _04691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12625__CLK clknet_leaf_172_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11764__I0 _05825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09820_ _04648_ _00633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06396__A1 u2.mem\[153\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09751_ _04605_ u2.mem\[37\]\[12\] _04606_ _04607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06963_ _02440_ _02441_ _02421_ _02442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_132_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08702_ _03722_ _03939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09682_ _04556_ _00587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06148__A1 u2.mem\[189\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06894_ _02365_ _02372_ _02353_ _02373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06148__B2 u2.mem\[176\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08633_ _03820_ u2.mem\[12\]\[9\] _03890_ _03892_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08564_ _03826_ u2.mem\[10\]\[12\] _03851_ _03852_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12005__CLK clknet_2_3__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11819__I1 u2.mem\[188\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07515_ u2.mem\[14\]\[7\] _02890_ _02891_ u2.mem\[12\]\[7\] _02987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07648__A1 u2.mem\[58\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08495_ _03807_ _00149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07446_ _02626_ _02920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08028__I _03488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06320__A1 u2.mem\[187\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06320__B2 u2.mem\[192\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10494__S _05061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07377_ u2.mem\[18\]\[4\] _02850_ _02851_ u2.mem\[19\]\[4\] _02852_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13400__CLK clknet_leaf_301_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09116_ _04132_ u2.mem\[23\]\[2\] _04203_ _04206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06328_ u2.mem\[152\]\[3\] _01712_ _01714_ u2.mem\[148\]\[3\] _01832_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08073__A1 _03523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09047_ _04160_ _04161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06259_ _01761_ _01762_ _01763_ _01764_ _01765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_135_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10007__I0 _04681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_83_clock_I clknet_5_9_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06387__A1 u2.mem\[158\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06387__B2 u2.mem\[151\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09949_ _04718_ _04729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_4002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11507__I0 _05680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12960_ _00839_ clknet_leaf_156_clock u2.mem\[52\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_1505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09523__S _04458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06011__I _01503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11911_ _03535_ _05929_ _05948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12891_ _00770_ clknet_leaf_219_clock u2.mem\[48\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_321_clock clknet_5_18_0_clock clknet_leaf_321_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07887__B2 u2.mem\[63\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11842_ _05903_ u2.mem\[190\]\[0\] _05905_ _05906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09322__I _04333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08687__I0 _03928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11773_ _05862_ _01372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13512_ _01391_ clknet_leaf_330_clock u2.mem\[188\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10494__I0 _05016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10724_ _05000_ _05204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06311__A1 u2.mem\[155\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_336_clock clknet_5_4_0_clock clknet_leaf_336_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13443_ _01322_ clknet_leaf_356_clock u2.mem\[177\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13080__CLK clknet_leaf_43_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10655_ _05112_ u2.mem\[59\]\[8\] _05162_ _05163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_360_clock_I clknet_5_0_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12648__CLK clknet_leaf_114_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13374_ _01253_ clknet_leaf_355_clock u2.mem\[165\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10586_ _05094_ _05122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_126_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12325_ _00204_ clknet_leaf_85_clock u2.mem\[12\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12256_ _00135_ clknet_leaf_228_clock u2.mem\[8\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11207_ _05508_ u2.mem\[150\]\[2\] _05502_ _05509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12798__CLK clknet_leaf_220_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12187_ _00066_ clknet_leaf_251_clock u2.mem\[4\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07575__B1 _02888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06378__B2 u2.mem\[155\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_11_0_clock_I clknet_3_5_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11138_ _05464_ u2.mem\[146\]\[1\] _05462_ _05465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08401__I _03484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12070__D data_in_trans\[10\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11069_ _04394_ _05402_ _05421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__12028__CLK clknet_leaf_307_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07017__I _02430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07878__A1 u2.mem\[53\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11426__A2 _05645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07300_ u2.mem\[8\]\[3\] _02612_ _02614_ u2.mem\[4\]\[3\] _02776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13423__CLK clknet_leaf_348_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10485__I0 _05007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08280_ _03659_ _03660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_32_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06302__A1 _01780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07231_ u2.mem\[58\]\[2\] _02495_ _02500_ u2.mem\[36\]\[2\] _02708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06853__A2 _02155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11203__S _05502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06591__I _02075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07162_ u2.mem\[15\]\[1\] _02457_ _02461_ u2.mem\[13\]\[1\] _02640_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13573__CLK clknet_leaf_20_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_105_clock_I clknet_5_11_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06113_ _01619_ _01607_ _01620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07093_ _02451_ _02452_ _02493_ _02544_ _02572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA_clkbuf_4_8_0_clock_I clknet_3_4_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08850__I0 _04030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09608__S _04511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06044_ col_select_trans\[4\].data_sync _01551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11737__I0 _05829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06369__A1 u2.mem\[146\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06369__B2 u2.mem\[186\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09407__I _04173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09803_ _04638_ _04639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06908__A3 _02353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08311__I _03684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06032__S _01510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07995_ _01562_ _01575_ _03458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_101_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09734_ _04592_ u2.mem\[37\]\[8\] _04593_ _04594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06946_ _02378_ _02421_ _02424_ _02425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_132_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09343__S _04346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07869__A1 u2.mem\[27\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09665_ _04469_ u2.mem\[36\]\[2\] _04544_ _04547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06877_ _02352_ _02353_ _02355_ _02356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08616_ _03882_ _00195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09596_ _04507_ _00550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08547_ _03842_ _00166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07090__C _02568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10476__I0 _04995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07097__A2 _02573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08478_ _03719_ u2.mem\[8\]\[14\] _03793_ _03796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07429_ u2.mem\[37\]\[5\] _02825_ _02826_ u2.mem\[59\]\[5\] _02903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06844__A2 _02114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10228__I0 _04898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08046__A1 _03503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10440_ _05033_ _00868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11976__I0 _05218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08841__I0 _04023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10371_ _04984_ _00848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12940__CLK clknet_leaf_256_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12110_ _05992_ clknet_leaf_18_clock u2.driver_enable vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09518__S _04453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13090_ _00969_ clknet_leaf_242_clock u2.mem\[60\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11728__I0 _05835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11847__I _03666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12041_ net3 clknet_2_3__leaf_clock_a col_select_trans\[2\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10751__I _05195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_307_clock_I clknet_5_16_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06780__A1 u2.mem\[155\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_260_clock clknet_5_23_0_clock clknet_leaf_260_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09253__S _04290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12943_ _00822_ clknet_leaf_237_clock u2.mem\[51\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10399__S _05002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12320__CLK clknet_leaf_158_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13446__CLK clknet_leaf_350_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12874_ _00753_ clknet_leaf_137_clock u2.mem\[46\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11825_ _05411_ _05886_ _05895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_2474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_275_clock clknet_5_21_0_clock clknet_leaf_275_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11756_ _05833_ u2.mem\[184\]\[3\] _05849_ _05853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12470__CLK clknet_leaf_106_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08824__A3 _03544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06296__B1 _01689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10707_ _05192_ _00976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06835__A2 _02100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11687_ _05786_ u2.mem\[180\]\[0\] _05810_ _05811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13426_ _01305_ clknet_leaf_349_clock u2.mem\[174\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10638_ _05153_ _00946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11967__I0 _05209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12065__D net21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11958__S _05975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13357_ _01236_ clknet_leaf_356_clock u2.mem\[163\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10862__S _05287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10569_ _03687_ _05110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06599__A1 _02023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_4_clock clknet_5_0_0_clock clknet_leaf_4_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12308_ _00187_ clknet_leaf_100_clock u2.mem\[11\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07260__A2 _02361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13288_ _01167_ clknet_leaf_364_clock u2.mem\[151\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_213_clock clknet_5_29_0_clock clknet_leaf_213_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_5_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11719__I0 _05829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12239_ _00118_ clknet_leaf_217_clock u2.mem\[7\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09227__I _04163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08131__I _03521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06800_ _02278_ _02279_ _02280_ _02281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07780_ u2.mem\[45\]\[12\] _03099_ _03100_ u2.mem\[34\]\[12\] _03247_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_228_clock clknet_5_25_0_clock clknet_leaf_228_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_83_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06771__A1 u2.mem\[171\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06771__B2 u2.mem\[157\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput4 col_select_a[3] net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06731_ _02210_ _02211_ _02212_ _02213_ _02214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_36_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09450_ _04391_ u2.mem\[30\]\[15\] _04411_ _04415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09560__I1 u2.mem\[33\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06662_ _02022_ _02012_ _02147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07720__B1 _03070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_31_clock_I clknet_5_3_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08401_ _03484_ _03749_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12813__CLK clknet_leaf_201_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09381_ _04147_ _04371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06593_ _02031_ _02077_ _02078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08332_ _03701_ _03702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06287__B1 _01734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08263_ _03648_ _00076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12963__CLK clknet_leaf_109_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07214_ u2.mem\[6\]\[1\] _02622_ _02624_ u2.mem\[47\]\[1\] _02692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08306__I _03680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08194_ _03482_ _03606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_118_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11958__I0 _05909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07145_ _02623_ _02624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_256_clock_I clknet_5_23_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13319__CLK clknet_leaf_301_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07251__A2 _02601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07076_ _02398_ _02399_ _02400_ _02552_ _02555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__08242__S _03635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06027_ u2.driver_mem\[14\] _01513_ _01535_ _01536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07003__A2 _02472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08041__I _03499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07085__C _02544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06211__B1 _01701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07978_ u2.mem\[26\]\[15\] _02573_ _02575_ u2.mem\[10\]\[15\] _03442_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_75_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06762__B2 u2.mem\[161\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09717_ _04579_ u2.mem\[37\]\[4\] _04580_ _04581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06929_ _02389_ _02408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_56_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11108__S _05445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10697__I0 _05117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09648_ _04536_ _00573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09579_ _04496_ u2.mem\[33\]\[14\] _04492_ _04497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11610_ _05750_ u2.mem\[175\]\[1\] _05761_ _05763_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12590_ _00469_ clknet_leaf_190_clock u2.mem\[29\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11110__I1 u2.mem\[144\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11541_ _05719_ u2.mem\[170\]\[5\] _05708_ _05720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11472_ _03506_ _05676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13211_ _01090_ clknet_leaf_287_clock u2.mem\[138\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10423_ _05022_ _00862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08814__I0 _03932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13142_ _01021_ clknet_leaf_23_clock u2.mem\[63\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10354_ _04902_ u2.mem\[52\]\[7\] _04971_ _04975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07242__A2 _02554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13073_ _00952_ clknet_leaf_236_clock u2.mem\[59\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10285_ _04935_ _00811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09047__I _04160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11177__I1 u2.mem\[148\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12024_ mem_address_trans\[9\].A clknet_leaf_289_clock mem_address_trans\[9\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08742__A2 _03606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12836__CLK clknet_leaf_61_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10688__I0 _05108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12926_ _00805_ clknet_leaf_255_clock u2.mem\[50\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07702__B1 _03112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12857_ _00736_ clknet_leaf_133_clock u2.mem\[45\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12986__CLK clknet_leaf_326_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11808_ _05876_ u2.mem\[187\]\[5\] _05878_ _05885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12788_ _00667_ clknet_leaf_71_clock u2.mem\[41\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11739_ _05831_ u2.mem\[183\]\[2\] _05840_ _05843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06808__A2 _02030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10860__I0 _05198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07481__A2 _02906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07030__I _02508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08805__I0 _03923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13409_ _01288_ clknet_leaf_305_clock u2.mem\[171\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07769__B1 _03081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_152_clock clknet_5_25_0_clock clknet_leaf_152_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_115_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07233__A2 _02654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12366__CLK clknet_leaf_209_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08950_ _04046_ u2.mem\[19\]\[14\] _04089_ _04092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07901_ _03363_ _03364_ _03365_ _03366_ _03367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08881_ _04052_ _00290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_167_clock clknet_5_26_0_clock clknet_leaf_167_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_69_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07832_ _02564_ _03299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09930__A1 _04288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06744__A1 u2.mem\[194\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06744__B2 u2.mem\[190\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07763_ u2.mem\[29\]\[11\] _03066_ _03067_ u2.mem\[11\]\[11\] _03231_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09502_ _04364_ u2.mem\[32\]\[3\] _04443_ _04447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06714_ _02133_ _02198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10679__I0 _05099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07694_ u2.mem\[40\]\[10\] _03018_ _03019_ u2.mem\[30\]\[10\] _03163_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09433_ _04405_ _00489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06645_ _02108_ _02070_ _02130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10767__S _05232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_09364_ _04359_ _00466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09297__I0 _04263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06576_ _02058_ _02053_ _02061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_105_clock clknet_5_11_0_clock clknet_leaf_105_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08315_ _03687_ _03688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10566__I _03683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09295_ _04260_ u2.mem\[27\]\[4\] _04318_ _04319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08246_ _03552_ u2.mem\[4\]\[3\] _03635_ _03639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10851__I0 _05204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07472__A2 _02893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08036__I data_in_trans\[1\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06275__A3 _01777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11598__S _05748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06680__B1 _02144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08177_ _03596_ _00042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12709__CLK clknet_leaf_27_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07128_ _02466_ _02467_ _02434_ _02483_ _02607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_134_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10007__S _04762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07059_ _02374_ _02538_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__13291__CLK clknet_leaf_361_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10070_ _04783_ _04802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12859__CLK clknet_leaf_199_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08700__S _03933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06735__A1 _02215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10972_ _05361_ _01072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12711_ _00590_ clknet_leaf_48_clock u2.mem\[36\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10677__S _05174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07160__A1 u2.mem\[27\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12642_ _00521_ clknet_leaf_174_clock u2.mem\[32\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09288__I0 _04254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06954__I _02432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12239__CLK clknet_leaf_217_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12573_ _00452_ clknet_leaf_187_clock u2.mem\[28\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11524_ _04287_ _05690_ _05708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_32_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12389__CLK clknet_leaf_78_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11455_ _05662_ _05663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_165_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07785__I _02414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11301__S _05568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10406_ _05010_ _00857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09460__I0 _04362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11386_ _05620_ _01227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13125_ _01004_ clknet_leaf_23_clock u2.mem\[62\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10337_ _04095_ _04964_ _04965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xclkbuf_leaf_84_clock clknet_5_11_0_clock clknet_leaf_84_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06974__A1 _02441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13056_ _00935_ clknet_leaf_243_clock u2.mem\[58\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09212__I0 _04265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10268_ _04891_ u2.mem\[50\]\[2\] _04923_ _04926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12007_ net25 clknet_2_2__leaf_clock_a mem_address_trans\[1\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10199_ _04879_ _00781_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_99_clock clknet_5_10_0_clock clknet_leaf_99_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11570__I1 u2.mem\[172\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_204_clock_I clknet_5_29_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13014__CLK clknet_leaf_28_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11971__S _05980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09441__S _04406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12909_ _00788_ clknet_leaf_202_clock u2.mem\[49\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_22_clock clknet_5_2_0_clock clknet_leaf_22_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07151__B2 u2.mem\[38\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06430_ u2.mem\[193\]\[1\] _01928_ _01929_ u2.mem\[192\]\[1\] _01914_ _01930_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_2090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09240__I _04176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13164__CLK clknet_leaf_270_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11086__I0 _05432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06361_ u2.mem\[153\]\[4\] _01708_ _01710_ u2.mem\[160\]\[4\] _01864_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08100_ _03481_ _03543_ _03544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xclkbuf_leaf_37_clock clknet_5_6_0_clock clknet_leaf_37_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_72_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09080_ _04185_ _00356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06292_ _01794_ _01795_ _01796_ _01797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08651__A1 _03901_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08031_ _03491_ _03492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput40 row_select_a[3] net40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11211__S _05502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11389__I1 u2.mem\[161\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07206__A2 _02601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10210__A1 _04013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09982_ _04696_ u2.mem\[43\]\[6\] _04745_ _04748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08933_ _04082_ _00312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06104__I _01610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08520__S _03818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11010__I0 _05384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08864_ _04040_ _00285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06717__A1 u2.mem\[194\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06717__B2 u2.mem\[190\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07815_ _02514_ _03282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08795_ _03989_ _03995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_45_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07390__A1 _02831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06193__A2 _01596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07746_ u2.mem\[50\]\[11\] _03111_ _03112_ u2.mem\[51\]\[11\] _03214_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_77_1100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13507__CLK clknet_leaf_330_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07677_ _02597_ _03147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09416_ _04395_ _04396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_129_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06628_ _02083_ _02090_ _02095_ _02112_ _02113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_129_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09150__I _04225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11077__I0 _05426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09347_ _04274_ u2.mem\[28\]\[10\] _04346_ _04349_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06559_ _02022_ _02044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12531__CLK clknet_leaf_103_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11777__A1 _04287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09278_ _04283_ u2.mem\[26\]\[14\] _04305_ _04308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09690__I0 _04494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08229_ _03577_ u2.mem\[3\]\[14\] _03624_ _03627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06653__B1 _02137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_0_clock_I clknet_5_0_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11240_ _05505_ u2.mem\[152\]\[1\] _05529_ _05531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12681__CLK clknet_leaf_129_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_153_clock_I clknet_5_25_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11171_ _05464_ u2.mem\[148\]\[1\] _05484_ _05486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06956__A1 _02429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10122_ _04834_ _00749_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13037__CLK clknet_leaf_267_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10053_ _04575_ _04790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06971__A4 _02449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06949__I _02427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06184__A2 _01615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11791__S _05865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12061__CLK clknet_2_0__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13187__CLK clknet_leaf_274_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_13_0_clock clknet_4_6_0_clock clknet_5_13_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_10955_ _05350_ _01066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_78_clock_I clknet_5_8_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10886_ _05305_ u2.mem\[130\]\[4\] _05296_ _05306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09060__I _04170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12625_ _00504_ clknet_leaf_172_clock u2.mem\[31\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09995__I _04739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12556_ _00435_ clknet_leaf_190_clock u2.mem\[27\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08605__S _03872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09681__I0 _04485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11507_ _05680_ u2.mem\[168\]\[5\] _05691_ _05698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07987__A3 _03449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10934__I _04117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12487_ _00366_ clknet_leaf_121_clock u2.mem\[22\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05998__A2 row_col_select_trans.data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11438_ _05635_ u2.mem\[164\]\[5\] _05646_ _05653_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12073__D net10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11369_ _05589_ u2.mem\[160\]\[2\] _05608_ _05611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11791__I1 u2.mem\[186\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13108_ _00987_ clknet_leaf_20_clock u2.mem\[61\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13039_ _00918_ clknet_leaf_320_clock u2.mem\[57\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09361__A2 _04250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_355_clock_I clknet_5_1_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07600_ u2.mem\[9\]\[8\] _03069_ _03070_ u2.mem\[25\]\[8\] _03071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08580_ _03806_ u2.mem\[11\]\[3\] _03857_ _03861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09171__S _04236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07531_ u2.mem\[17\]\[7\] _02844_ _02845_ u2.mem\[24\]\[7\] _03003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12554__CLK clknet_leaf_119_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10110__S _04825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07462_ u2.mem\[16\]\[6\] _02798_ _02799_ u2.mem\[33\]\[6\] _02935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06594__I _02078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09201_ _04135_ _04258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06413_ _01913_ _01914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07393_ _02447_ _02867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09132_ _04158_ u2.mem\[23\]\[9\] _04213_ _04215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06344_ u2.mem\[172\]\[4\] _01654_ _01667_ u2.mem\[150\]\[4\] _01847_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07427__A2 _02899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09672__I0 _04476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09063_ data_in_trans\[14\].data_sync _04173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07639__B _02978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06275_ _01771_ _01774_ _01777_ _01779_ _01780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_135_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08014_ u3.enable _03476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08314__I data_in_trans\[7\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11231__I0 _05514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10780__S _05237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09965_ _04716_ u2.mem\[42\]\[15\] _04734_ _04738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08916_ _04071_ _04072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_4206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12084__CLK clknet_leaf_363_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09896_ _04694_ u2.mem\[41\]\[5\] _04692_ _04695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08847_ _04028_ u2.mem\[17\]\[6\] _04024_ _04029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07093__C _02544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07363__A1 u2.mem\[9\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07363__B2 u2.mem\[25\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08984__I _04096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08778_ _03982_ _00257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09081__S _04182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07729_ u2.mem\[39\]\[10\] _03088_ _03089_ u2.mem\[48\]\[10\] _03198_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_1553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10020__S _04767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10740_ _05215_ _00986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_5_31_0_clock_I clknet_4_15_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10671_ _05171_ _00961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12410_ _00289_ clknet_leaf_112_clock u2.mem\[17\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07418__A2 _02890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13390_ _01269_ clknet_leaf_355_clock u2.mem\[168\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06009__I _01507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09663__I0 _04467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12341_ _00220_ clknet_leaf_79_clock u2.mem\[13\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11470__I0 _05674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10754__I _03713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12272_ _00151_ clknet_leaf_166_clock u2.mem\[9\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08224__I _03608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11223_ _05500_ u2.mem\[151\]\[0\] _05520_ _05521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10690__S _05179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09256__S _04295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08160__S _03585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11154_ _05460_ u2.mem\[147\]\[0\] _05475_ _05476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10105_ _04819_ _04825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_1_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11085_ _05351_ _05432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09055__I _04166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10036_ _04712_ u2.mem\[44\]\[13\] _04777_ _04779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12577__CLK clknet_leaf_170_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11987_ _01979_ _05972_ _05991_ _01457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11026__S _05395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10938_ _05335_ u2.mem\[134\]\[0\] _05337_ _05338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07121__A4 _02498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12068__D data_in_trans\[9\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10869_ _05293_ _01037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12608_ _00487_ clknet_leaf_172_clock u2.mem\[30\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07409__A2 _02881_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09654__I0 _04496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12539_ _00418_ clknet_leaf_184_clock u2.mem\[26\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13202__CLK clknet_leaf_280_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07290__B1 _02582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08134__I _03523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06060_ _01566_ _01567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11913__A1 _04013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11764__I1 u2.mem\[185\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13352__CLK clknet_leaf_361_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07593__A1 _03054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06396__A2 _01707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06962_ _02409_ _02441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09750_ _04566_ _04606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_136_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08701_ _03938_ _00224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09681_ _04485_ u2.mem\[36\]\[9\] _04554_ _04556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06893_ _02339_ _02338_ _02344_ _02372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07345__A1 _02791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08632_ _03891_ _00202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_101_clock_I clknet_5_11_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08563_ _03835_ _03851_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_81_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08145__I0 _03575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07514_ u2.mem\[44\]\[7\] _02887_ _02888_ u2.mem\[42\]\[7\] _02986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08494_ _03806_ u2.mem\[9\]\[3\] _03800_ _03807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08309__I data_in_trans\[6\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09893__I0 _04691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07445_ _02915_ _02916_ _02917_ _02918_ _02919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_126_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06320__A2 _01632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07376_ _02607_ _02851_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09645__I0 _04487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09115_ _04205_ _00371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11452__I0 _05635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06327_ u2.mem\[153\]\[3\] _01707_ _01709_ u2.mem\[160\]\[3\] _01831_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08073__A2 _03519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09046_ data_in_trans\[10\].data_sync _04160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08044__I data_in_trans\[3\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06258_ u2.mem\[189\]\[1\] _01649_ _01651_ u2.mem\[176\]\[1\] u2.mem\[172\]\[1\]
+ _01653_ _01764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_136_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07820__A2 _03132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_26_clock_I clknet_5_2_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06189_ _01685_ _01690_ _01695_ _01696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_46_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07033__B1 _02511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06926__A4 _02404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06499__I row_select_trans\[0\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09948_ _04728_ _00681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11507__I1 u2.mem\[168\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06792__C1 u2.mem\[168\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09804__S _04639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07336__A1 u2.mem\[58\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09879_ _04682_ _04683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_4047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11910_ _05947_ _01424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12890_ _00769_ clknet_leaf_140_clock u2.mem\[47\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07887__A2 _02559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09603__I _04500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10891__A1 _04072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11841_ _05904_ _05905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_166_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07639__A2 _03034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11772_ _05835_ u2.mem\[185\]\[4\] _05856_ _05862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06847__B1 _02130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13511_ _01390_ clknet_leaf_317_clock u2.mem\[188\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10723_ _05203_ _00981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11691__I0 _05792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10494__I1 u2.mem\[55\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13225__CLK clknet_leaf_283_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13442_ _01321_ clknet_leaf_356_clock u2.mem\[177\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10654_ _05151_ _05162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_139_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09636__I0 _04478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_303_clock_I clknet_5_16_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13373_ _01252_ clknet_leaf_354_clock u2.mem\[165\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10585_ _03708_ _05121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12324_ _00203_ clknet_leaf_84_clock u2.mem\[12\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07272__B1 _02646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07811__A2 _03271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12255_ _00134_ clknet_leaf_217_clock u2.mem\[8\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11206_ _05507_ _05508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12186_ _00065_ clknet_leaf_59_clock u2.mem\[3\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11137_ _05339_ _05464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11068_ _05334_ _05420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10019_ _04769_ _00711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_4_15_0_clock_I clknet_3_7_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09513__I _04442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09875__I0 _04615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11682__I0 _05798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06302__A2 _01784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07230_ u2.mem\[53\]\[2\] _02486_ _02489_ u2.mem\[56\]\[2\] _02707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09627__I0 _04469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07161_ _02635_ _02636_ _02637_ _02638_ _02639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__11434__I0 _05631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10394__I _04988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06112_ _01558_ _01568_ _01585_ _01619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_146_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07092_ u2.mem\[29\]\[0\] _02565_ _02570_ u2.mem\[11\]\[0\] _02571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06043_ col_select_trans\[5\].data_sync _01550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07917__B _03211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12742__CLK clknet_leaf_70_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11737__I1 u2.mem\[183\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06369__A2 _01691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09802_ _03752_ _04542_ _04638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_140_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07994_ _01980_ _03246_ _03436_ _03457_ _01492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12892__CLK clknet_leaf_209_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09733_ _04566_ _04593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06945_ _02349_ _02423_ _02424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_132_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07581__A4 _03051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09664_ _04546_ _00579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06876_ _02339_ _02354_ _02355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_252_clock_I clknet_5_22_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08615_ _03802_ u2.mem\[12\]\[1\] _03880_ _03882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09595_ _04473_ u2.mem\[34\]\[4\] _04506_ _04507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10569__I _03687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12122__CLK clknet_leaf_328_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13248__CLK clknet_leaf_272_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08546_ _03808_ u2.mem\[10\]\[4\] _03841_ _03842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09866__I0 _04602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08477_ _03795_ _00143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07428_ u2.mem\[60\]\[5\] _02822_ _02823_ u2.mem\[62\]\[5\] _02902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12272__CLK clknet_leaf_166_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13398__CLK clknet_leaf_307_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07359_ _02569_ _02834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07254__B1 _02688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10370_ _04918_ u2.mem\[52\]\[14\] _04981_ _04984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08703__S _03933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09029_ data_in_trans\[6\].data_sync _04147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12040_ col_select_trans\[1\].A clknet_leaf_299_clock col_select_trans\[1\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09534__S _04465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07309__A1 u2.mem\[32\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06780__A2 _02029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06957__I _02435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12942_ _00821_ clknet_leaf_255_clock u2.mem\[51\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09333__I _04335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12873_ _00752_ clknet_leaf_137_clock u2.mem\[46\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08109__I0 _03550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11824_ _05894_ _01391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09857__I0 _04589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12615__CLK clknet_leaf_113_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11755_ _05852_ _01364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07788__I _02435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06296__A1 u2.mem\[170\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06296__B2 u2.mem\[156\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10706_ _05126_ u2.mem\[60\]\[14\] _05189_ _05192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11686_ _05809_ _05810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_13425_ _01304_ clknet_leaf_349_clock u2.mem\[174\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10637_ _05093_ u2.mem\[59\]\[0\] _05152_ _05153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11103__I _05442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07245__B1 _02570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08613__S _03880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13356_ _01235_ clknet_leaf_360_clock u2.mem\[162\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10568_ _05109_ _00920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06599__A2 _02058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07796__B2 u2.mem\[7\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12307_ _00186_ clknet_leaf_104_clock u2.mem\[11\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13287_ _01166_ clknet_leaf_364_clock u2.mem\[151\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10499_ _05020_ u2.mem\[55\]\[12\] _05066_ _05067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11719__I1 u2.mem\[182\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12238_ _00117_ clknet_leaf_211_clock u2.mem\[7\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08596__I0 _03822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12081__D net45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12169_ _00048_ clknet_leaf_131_clock u2.mem\[2\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12145__CLK clknet_leaf_218_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06771__A2 _02065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06730_ u2.mem\[180\]\[2\] _02043_ _02014_ u2.mem\[172\]\[2\] _02213_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput5 col_select_a[4] net5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06661_ _02145_ _02146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10389__I _04997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07720__B2 u2.mem\[25\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08400_ _03605_ _03482_ _03748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09380_ _04370_ _00471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12295__CLK clknet_leaf_120_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06592_ _02026_ _01991_ _02077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09848__I0 _04576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08331_ _03700_ _03701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13540__CLK clknet_leaf_34_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08520__I0 _03824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06287__A1 u2.mem\[193\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08262_ _03568_ u2.mem\[4\]\[10\] _03645_ _03648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06287__B2 u2.mem\[177\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07213_ u2.mem\[8\]\[1\] _02612_ _02614_ u2.mem\[4\]\[1\] _02691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08193_ mem_address_trans\[1\].data_sync _03605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_146_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06039__A1 col_select_trans\[0\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07236__B1 _02517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07144_ _02469_ _02491_ _02492_ _02453_ _02623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_9_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11958__I1 u2.mem\[194\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_320_clock clknet_5_18_0_clock clknet_leaf_320_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_160_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07075_ _02553_ _02554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06026_ u2.driver_mem\[15\] _01508_ _01535_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_126_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08322__I _03659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08587__I0 _03813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_335_clock clknet_5_5_0_clock clknet_leaf_335_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_102_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input37_I row_select_a[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06211__A1 u2.mem\[154\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06211__B2 u2.mem\[162\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07977_ _03437_ _03438_ _03439_ _03440_ _03441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_56_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13070__CLK clknet_leaf_253_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09716_ _04566_ _04580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_132_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06928_ _02387_ _02407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_67_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12638__CLK clknet_leaf_192_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09647_ _04489_ u2.mem\[35\]\[11\] _04532_ _04536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06859_ _02009_ row_select_trans\[4\].data_sync _02338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_56_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09578_ _04173_ _04496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08529_ _03718_ _03831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11646__I0 _05756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12788__CLK clknet_leaf_71_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08511__I0 _03817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11124__S _05453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06278__B2 u2.mem\[150\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11540_ _05679_ _05719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11471_ _05675_ _01257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10963__S _05356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09529__S _04458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12018__CLK clknet_leaf_299_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13210_ _01089_ clknet_leaf_281_clock u2.mem\[138\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10422_ _05020_ u2.mem\[53\]\[12\] _05021_ _05022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07778__A1 _01966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10353_ _04974_ _00840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13141_ _01020_ clknet_leaf_19_clock u2.mem\[63\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13072_ _00951_ clknet_leaf_241_clock u2.mem\[59\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10284_ _04907_ u2.mem\[50\]\[9\] _04933_ _04935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08578__I0 _03804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12168__CLK clknet_leaf_109_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12023_ net33 clknet_2_1__leaf_clock_a mem_address_trans\[9\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11794__S _05865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13413__CLK clknet_leaf_344_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06202__A1 _01600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07950__A1 _03399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10203__S _04880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09063__I data_in_trans\[14\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13563__CLK clknet_leaf_16_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12925_ _00804_ clknet_leaf_257_clock u2.mem\[50\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11885__I0 u2.mem\[192\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08750__I0 _03912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_148_clock_I clknet_5_24_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12856_ _00735_ clknet_leaf_129_clock u2.mem\[45\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11807_ _05884_ _01384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10937__I _05336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12787_ _00666_ clknet_leaf_26_clock u2.mem\[41\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11034__S _05394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06269__A1 u2.mem\[178\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06269__B2 u2.mem\[164\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07466__B1 _02882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11738_ _05842_ _01357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07311__I _02414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11969__S _05980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12076__D data_in_trans\[13\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11669_ _05799_ _01331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_200_clock_I clknet_5_28_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09439__S _04406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07218__B1 _02634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13408_ _01287_ clknet_leaf_304_clock u2.mem\[171\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10672__I _04862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13339_ _01218_ clknet_leaf_4_clock u2.mem\[160\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07900_ u2.mem\[18\]\[13\] _03316_ _03317_ u2.mem\[19\]\[13\] _03366_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13093__CLK clknet_leaf_24_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08880_ _04010_ u2.mem\[18\]\[0\] _04051_ _04052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07831_ u2.mem\[26\]\[12\] _03139_ _03140_ u2.mem\[10\]\[12\] _03298_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09930__A2 _04659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06597__I _02081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07762_ u2.mem\[26\]\[11\] _03139_ _03140_ u2.mem\[10\]\[11\] _03230_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10128__I0 _04815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09501_ _04446_ _00516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06713_ u2.mem\[153\]\[1\] _02196_ _02131_ u2.mem\[152\]\[1\] _02197_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07693_ u2.mem\[32\]\[10\] _03015_ _03016_ u2.mem\[2\]\[10\] _03162_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09432_ _04373_ u2.mem\[30\]\[7\] _04401_ _04405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06644_ _02128_ _02129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11628__I0 _05752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09363_ _04356_ u2.mem\[29\]\[0\] _04358_ _04359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06575_ _02059_ _02060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09297__I1 u2.mem\[27\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08314_ data_in_trans\[7\].data_sync _03687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09294_ _04312_ _04318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_123_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08245_ _03638_ _00068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10783__S _05242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09349__S _04346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11005__A1 _04288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08176_ _03563_ u2.mem\[2\]\[8\] _03595_ _03596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06680__B2 u2.mem\[147\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07127_ _02605_ _02606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11800__I0 _05868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13436__CLK clknet_leaf_350_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09148__I _04223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07058_ _02370_ _02537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_161_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06983__A2 _02457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_274_clock clknet_5_21_0_clock clknet_leaf_274_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06009_ _01507_ _01518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12460__CLK clknet_leaf_196_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08980__I0 _04037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10119__I0 _04806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_289_clock clknet_5_20_0_clock clknet_leaf_289_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_29_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11867__I0 _05911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10971_ _05349_ u2.mem\[135\]\[4\] _05355_ _05361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10958__S _05336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12710_ _00589_ clknet_leaf_27_clock u2.mem\[36\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_3_clock clknet_5_0_0_clock clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07160__A2 _02428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_212_clock clknet_5_29_0_clock clknet_leaf_212_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12641_ _00520_ clknet_leaf_173_clock u2.mem\[32\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10757__I _03717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09288__I1 u2.mem\[27\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07448__B1 _02921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12572_ _00451_ clknet_leaf_186_clock u2.mem\[28\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11523_ _05662_ _05707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10693__S _05184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_227_clock clknet_5_25_0_clock clknet_leaf_227_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_172_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11454_ _03491_ _05662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11588__I _05747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10405_ _05009_ u2.mem\[53\]\[7\] _05002_ _05010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11385_ _05591_ u2.mem\[161\]\[3\] _05616_ _05620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09460__I1 u2.mem\[31\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13124_ _01003_ clknet_leaf_23_clock u2.mem\[62\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10336_ _04862_ _04964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12803__CLK clknet_leaf_145_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_74_clock_I clknet_5_8_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08897__I _04050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10267_ _04925_ _00803_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13055_ _00934_ clknet_leaf_240_clock u2.mem\[58\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12006_ mem_address_trans\[0\].A clknet_leaf_312_clock mem_address_trans\[0\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06411__S _01502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10198_ _04808_ u2.mem\[48\]\[11\] _04875_ _04879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07923__A1 _03384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06726__A2 _02206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08971__I0 _04028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12953__CLK clknet_leaf_324_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10868__S _05286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_299_clock_I clknet_5_17_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12908_ _00787_ clknet_leaf_202_clock u2.mem\[49\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07687__B1 _03092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08338__S _03694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10530__I0 _05014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07151__A2 _02627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13309__CLK clknet_leaf_348_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12839_ _00718_ clknet_leaf_135_clock u2.mem\[44\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06360_ u2.mem\[190\]\[4\] _01703_ _01705_ u2.mem\[194\]\[4\] _01863_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08137__I _03525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12333__CLK clknet_leaf_209_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06291_ u2.mem\[152\]\[2\] _01713_ _01715_ u2.mem\[148\]\[2\] _01796_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10833__I1 _03533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08030_ data_in_trans\[0\].data_sync _03491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09169__S _04236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06880__I _02358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06662__A1 _02022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput30 mem_address_a[6] net30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput41 row_select_a[4] net41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10108__S _04825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12483__CLK clknet_leaf_123_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07611__B1 _03081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10210__A2 _04863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09981_ _04747_ _00695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08954__A3 _03633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08932_ _04028_ u2.mem\[19\]\[6\] _04079_ _04082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08600__I _03856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08863_ _04039_ u2.mem\[17\]\[11\] _04033_ _04040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08962__I0 _04019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07814_ u2.mem\[49\]\[12\] _03126_ _03127_ u2.mem\[46\]\[12\] _03281_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08794_ _03994_ _00261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09632__S _04527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07390__A2 _02842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07745_ _03208_ _03209_ _03210_ _03212_ _03213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10778__S _05237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07678__B1 _03147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07676_ _02595_ _03146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10521__I0 _05005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09415_ _04394_ _04011_ _04395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_13_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06627_ u2.mem\[166\]\[0\] _02097_ _02099_ u2.mem\[161\]\[0\] _02111_ _02112_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_40_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09346_ _04348_ _00459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06558_ _02042_ _02043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11777__A2 _05847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10824__I1 _03523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09277_ _04307_ _00431_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06489_ u2.mem\[0\]\[14\] _01976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09690__I1 u2.mem\[36\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09079__S _04182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06653__A1 u2.mem\[153\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08228_ _03626_ _00063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06653__B2 u2.mem\[160\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12826__CLK clknet_leaf_136_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08159_ _03586_ _00034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10018__S _04767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11201__I _03496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11170_ _05485_ _01146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08711__S _03942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10121_ _04808_ u2.mem\[46\]\[11\] _04830_ _04834_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12976__CLK clknet_leaf_249_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10052_ _04789_ _00724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08510__I _03799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12206__CLK clknet_leaf_212_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10688__S _05179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06965__I _02443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_151_clock clknet_5_25_0_clock clknet_leaf_151_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08158__S _03585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10954_ _05349_ u2.mem\[134\]\[4\] _05336_ _05350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10512__I0 _04992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12356__CLK clknet_leaf_80_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10885_ _05000_ _05305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12624_ _00503_ clknet_leaf_168_clock u2.mem\[31\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09130__I0 _04154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_166_clock clknet_5_26_0_clock clknet_leaf_166_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_129_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12555_ _00434_ clknet_leaf_191_clock u2.mem\[27\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10815__I1 _03513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11506_ _05697_ _01270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12486_ _00365_ clknet_leaf_100_clock u2.mem\[22\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11437_ _05652_ _01246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11368_ _05610_ _01219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13107_ _00986_ clknet_leaf_20_clock u2.mem\[61\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10319_ _04904_ u2.mem\[51\]\[8\] _04954_ _04955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11299_ _04333_ _05566_ _05567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_80_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_104_clock clknet_5_11_0_clock clknet_leaf_104_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13038_ _00917_ clknet_leaf_248_clock u2.mem\[57\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11982__S _05985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07036__I _02514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11781__I _03662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_119_clock clknet_5_15_0_clock clknet_leaf_119_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_130_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07530_ u2.mem\[23\]\[7\] _02913_ _02914_ u2.mem\[22\]\[7\] _03002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11456__A1 _04179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10503__I0 _05025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07461_ u2.mem\[1\]\[6\] _02795_ _02796_ u2.mem\[7\]\[6\] _02934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10397__I _04143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06332__B1 _01689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13281__CLK clknet_leaf_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09200_ _04257_ _00404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06412_ _01911_ _01912_ _01913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06883__A1 _02338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07392_ _02443_ _02866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12849__CLK clknet_leaf_154_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09121__I0 _04140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09131_ _04214_ _00378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06343_ u2.mem\[174\]\[4\] _01657_ _01659_ u2.mem\[155\]\[4\] _01661_ u2.mem\[181\]\[4\]
+ _01846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__10806__I1 _03500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06824__B _02304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09062_ _04172_ _00351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06274_ u2.mem\[184\]\[2\] _01778_ _01554_ _01779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_159_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08013_ _03468_ _03475_ _05992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12999__CLK clknet_leaf_323_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11021__I _05351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09627__S _04522_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11231__I1 u2.mem\[151\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06399__B1 _01701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07060__A1 _02455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09964_ _04737_ _00688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12229__CLK clknet_leaf_69_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08915_ _03485_ _03748_ _04071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08330__I data_in_trans\[10\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09895_ _04582_ _04694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11892__S _05937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08846_ _03684_ _04028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10742__I0 _05216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08777_ _03939_ u2.mem\[15\]\[15\] _03978_ _03982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12379__CLK clknet_leaf_207_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07728_ u2.mem\[5\]\[10\] _03153_ _03154_ u2.mem\[38\]\[10\] _03197_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10301__S _04944_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07115__A2 _02591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_22_clock_I clknet_5_2_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07659_ u2.mem\[43\]\[9\] _03049_ _03050_ u2.mem\[20\]\[9\] _03129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_83_clock clknet_5_9_0_clock clknet_leaf_83_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_25_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10670_ _05128_ u2.mem\[59\]\[15\] _05167_ _05171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09112__I0 _04119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09329_ _04256_ u2.mem\[28\]\[2\] _04336_ _04339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09663__I1 u2.mem\[36\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12340_ _00219_ clknet_leaf_80_clock u2.mem\[13\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_98_clock clknet_5_10_0_clock clknet_leaf_98_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_126_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13004__CLK clknet_leaf_257_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12271_ _00150_ clknet_leaf_166_clock u2.mem\[9\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10971__S _05355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09537__S _04465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11222_ _05519_ _05520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_134_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_21_clock clknet_5_2_0_clock clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07051__A1 _02413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11153_ _05474_ _05475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_96_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10104_ _04824_ _00741_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13154__CLK clknet_leaf_263_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11084_ _05431_ _01114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10035_ _04778_ _00718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08000__B1 _03462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_36_clock clknet_5_4_0_clock clknet_leaf_36_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_76_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11307__S _05568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11986_ _03535_ _05972_ _05991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10937_ _05336_ _05337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_31_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10868_ _05207_ u2.mem\[129\]\[5\] _05286_ _05293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12607_ _00486_ clknet_leaf_173_clock u2.mem\[30\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10945__I _05342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_10799_ _05251_ _01009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06617__A1 u2.mem\[187\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12538_ _00417_ clknet_leaf_115_clock u2.mem\[25\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07814__B1 _03127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08415__I _03753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06617__B2 u2.mem\[192\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12469_ _00348_ clknet_leaf_106_clock u2.mem\[21\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11776__I _03655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11913__A2 _05926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09246__I _04289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08150__I _03535_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06961_ _02348_ _02423_ _02440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_08700_ _03937_ u2.mem\[13\]\[14\] _03933_ _03938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12521__CLK clknet_leaf_118_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09680_ _04555_ _00586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06892_ _02370_ _02371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_39_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09590__I0 _04469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08631_ _03817_ u2.mem\[12\]\[8\] _03890_ _03891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08562_ _03850_ _00173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10121__S _04830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07513_ _02981_ _02982_ _02983_ _02984_ _02985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA_clkbuf_leaf_196_clock_I clknet_5_31_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08493_ _03671_ _03806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09893__I1 u2.mem\[41\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07444_ u2.mem\[18\]\[5\] _02850_ _02851_ u2.mem\[19\]\[5\] _02918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07375_ _02605_ _02850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13027__CLK clknet_leaf_42_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09114_ _04128_ u2.mem\[23\]\[1\] _04203_ _04205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06608__A1 _02031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06326_ u2.mem\[190\]\[3\] _01702_ _01704_ u2.mem\[194\]\[3\] _01830_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08325__I data_in_trans\[9\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11452__I1 u2.mem\[165\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11887__S _05932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09045_ _04159_ _00347_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06257_ u2.mem\[190\]\[1\] _01703_ _01710_ u2.mem\[160\]\[1\] _01705_ u2.mem\[194\]\[1\]
+ _01763_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_50_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12051__CLK clknet_2_0__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13177__CLK clknet_leaf_275_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06188_ u2.mem\[146\]\[0\] _01692_ _01694_ u2.mem\[186\]\[0\] _01695_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11686__I _05809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10963__I0 _05335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09947_ _04698_ u2.mem\[42\]\[7\] _04724_ _04728_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06792__B1 _02086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06792__C2 _02093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08995__I _04118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09878_ _04249_ _04659_ _04682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08829_ _04016_ _00274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10031__S _04772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11840_ _04393_ _05886_ _05904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_2635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07404__I _02502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06448__C _01934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11771_ _05861_ _01371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13510_ _01389_ clknet_leaf_335_clock u2.mem\[188\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10722_ _05202_ u2.mem\[61\]\[3\] _05196_ _05203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08436__S _03769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06847__B2 u2.mem\[152\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11840__A1 _04393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11691__I1 u2.mem\[180\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13441_ _01320_ clknet_leaf_348_clock u2.mem\[177\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10653_ _05161_ _00953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13372_ _01251_ clknet_leaf_359_clock u2.mem\[165\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10584_ _05120_ _00925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12323_ _00202_ clknet_leaf_84_clock u2.mem\[12\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09267__S _04300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12254_ _00133_ clknet_leaf_216_clock u2.mem\[8\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11205_ _03499_ _05507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12544__CLK clknet_leaf_168_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12185_ _00064_ clknet_leaf_59_clock u2.mem\[3\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10954__I0 _05349_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07575__A2 _02887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11136_ _05463_ _01134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11067_ _05419_ _01109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10706__I0 _05126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10018_ _04694_ u2.mem\[44\]\[5\] _04767_ _04769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07314__I _02435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06358__C _01860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12079__D net13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11969_ _05211_ u2.mem\[194\]\[7\] _05980_ _05982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06302__A3 _01793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06374__B _01876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07160_ u2.mem\[27\]\[1\] _02428_ _02436_ u2.mem\[35\]\[1\] _02638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12074__CLK clknet_leaf_343_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11434__I1 u2.mem\[164\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06111_ _01615_ _01617_ _01618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_157_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07263__A1 u2.mem\[40\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07091_ _02569_ _02570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06042_ _01548_ _01549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07015__A1 _02413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09801_ _04637_ _00625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07993_ _03441_ _03446_ _03451_ _03456_ _03457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_140_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09732_ _04591_ _04592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_171_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06944_ _02422_ _02350_ _02423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09563__I0 _04485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09663_ _04467_ u2.mem\[36\]\[1\] _04544_ _04546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06875_ row_select_trans\[1\].data_sync _02010_ _02354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08614_ _03881_ _00194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09594_ _04500_ _04506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_43_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09315__I0 _04281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08545_ _03835_ _03841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_42_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11122__I0 _05424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09866__I1 u2.mem\[40\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12417__CLK clknet_leaf_161_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08476_ _03715_ u2.mem\[8\]\[13\] _03793_ _03795_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07427_ u2.mem\[61\]\[5\] _02899_ _02900_ u2.mem\[63\]\[5\] _02901_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10585__I _03708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08055__I _03510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07358_ _02564_ _02833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06309_ u2.mem\[184\]\[3\] _01778_ _01749_ _01813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12567__CLK clknet_leaf_113_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07254__B2 u2.mem\[38\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07289_ u2.mem\[29\]\[3\] _02565_ _02570_ u2.mem\[11\]\[3\] _02765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_152_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09028_ _04146_ _00343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11189__I0 _05468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07006__A1 _02483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12941_ _00820_ clknet_leaf_256_clock u2.mem\[51\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12872_ _00751_ clknet_leaf_137_clock u2.mem\[46\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07190__B1 _02667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09306__I0 _04272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09550__S _04474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11823_ _05876_ u2.mem\[188\]\[5\] _05887_ _05894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06973__I _02408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11754_ _05831_ u2.mem\[184\]\[2\] _05849_ _05852_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13342__CLK clknet_leaf_4_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10705_ _05191_ _00975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07493__A1 u2.mem\[8\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11685_ _04094_ _05808_ _05809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_122_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13424_ _01303_ clknet_leaf_347_clock u2.mem\[174\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10636_ _05151_ _05152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_167_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07245__A1 u2.mem\[29\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13355_ _01234_ clknet_leaf_360_clock u2.mem\[162\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13492__CLK clknet_leaf_292_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10567_ _05108_ u2.mem\[57\]\[6\] _05104_ _05109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12306_ _00185_ clknet_leaf_166_clock u2.mem\[11\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_144_clock_I clknet_5_24_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13286_ _01165_ clknet_leaf_1_clock u2.mem\[151\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10498_ _05050_ _05066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_29_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12237_ _00116_ clknet_leaf_211_clock u2.mem\[7\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06213__I _01719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12168_ _00047_ clknet_leaf_109_clock u2.mem\[2\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11119_ _05452_ _05453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_12099_ _01497_ clknet_leaf_149_clock u2.active_mem\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput6 col_select_a[5] net6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06660_ _02057_ _02125_ _02145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07181__B1 _02658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07720__A2 _03069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09460__S _04419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06591_ _02075_ _02076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09848__I1 u2.mem\[40\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_69_clock_I clknet_5_9_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08330_ data_in_trans\[10\].data_sync _03700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07079__A4 _02442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08261_ _03647_ _00075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07212_ u2.mem\[39\]\[1\] _02617_ _02619_ u2.mem\[48\]\[1\] _02690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_14_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08192_ _03604_ _00049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06039__A2 col_select_trans\[1\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07143_ _02621_ _02622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07236__B2 u2.mem\[20\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07074_ _02551_ _02537_ _02538_ _02552_ _02553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_12_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06025_ _01516_ _01533_ _01534_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10918__I0 _05307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08587__I1 u2.mem\[11\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13215__CLK clknet_leaf_283_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06211__A2 _01699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07976_ u2.mem\[57\]\[15\] _03294_ _03295_ u2.mem\[41\]\[15\] _03440_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_19_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09434__I _04395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09715_ _04578_ _04579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06927_ _02405_ _02406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_346_clock_I clknet_5_4_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09646_ _04535_ _00572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06858_ _01878_ _01996_ _02337_ _01479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11894__I1 _03515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07172__B1 _02649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13365__CLK clknet_leaf_358_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09577_ _04495_ _00543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06789_ _02255_ _02260_ _02265_ _02270_ _02271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08528_ _03830_ _00159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07475__A1 _02932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06278__A2 _01654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08459_ _03785_ _00135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11470_ _05674_ u2.mem\[166\]\[3\] _05665_ _05675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10421_ _04988_ _05021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07778__A2 _03013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13140_ _01019_ clknet_leaf_22_clock u2.mem\[63\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10352_ _04900_ u2.mem\[52\]\[6\] _04971_ _04974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08513__I _03697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13071_ _00950_ clknet_leaf_240_clock u2.mem\[59\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10283_ _04934_ _00810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07129__I _02607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12022_ mem_address_trans\[8\].A clknet_leaf_287_clock mem_address_trans\[8\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11582__I0 _05717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06202__A2 _01634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08742__A4 _03878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09527__I0 _04389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07950__A2 _03404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12924_ _00803_ clknet_leaf_257_clock u2.mem\[50\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07163__B1 _02471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11885__I1 _03503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09280__S _04305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07702__A2 _03111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12855_ _00734_ clknet_leaf_133_clock u2.mem\[45\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_70_clock_I clknet_5_8_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11315__S _05576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11806_ _05874_ u2.mem\[187\]\[4\] _05878_ _05884_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12786_ _00665_ clknet_leaf_321_clock u2.mem\[41\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11737_ _05829_ u2.mem\[183\]\[1\] _05840_ _05842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06208__I _01714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08624__S _03885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11668_ _05798_ u2.mem\[178\]\[5\] _05787_ _05799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12882__CLK clknet_leaf_230_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13407_ _01286_ clknet_leaf_304_clock u2.mem\[171\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10619_ _05142_ _00938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10953__I _05348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11599_ _05755_ _01305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07769__A2 _03080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13338_ _01217_ clknet_leaf_9_clock u2.mem\[159\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_295_clock_I clknet_5_17_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12092__D inverter_select_trans.A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13269_ _01148_ clknet_leaf_5_clock u2.mem\[148\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11784__I _03666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07830_ _03287_ _03290_ _03293_ _03296_ _03297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_57_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12262__CLK clknet_leaf_69_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09518__I0 _04380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13388__CLK clknet_leaf_355_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07761_ _03225_ _03226_ _03227_ _03228_ _03229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_42_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11325__I0 _05556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09500_ _04362_ u2.mem\[32\]\[2\] _04443_ _04446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06712_ _02136_ _02196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07692_ u2.mem\[45\]\[10\] _03099_ _03100_ u2.mem\[34\]\[10\] _03161_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09431_ _04404_ _00488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06643_ _02108_ _02041_ _02128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11225__S _05520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09362_ _04357_ _04358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11628__I1 u2.mem\[176\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06574_ _02057_ _02058_ _02059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08313_ _03686_ _00088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07457__A1 u2.mem\[40\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09293_ _04317_ _00437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08244_ _03550_ u2.mem\[4\]\[2\] _03635_ _03638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08175_ _03584_ _03595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_118_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06680__A2 _02142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10064__I0 _04797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07126_ _02566_ _02567_ _02393_ _02547_ _02605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_146_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11800__I1 u2.mem\[187\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07057_ _02450_ _02482_ _02513_ _02535_ _02536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_106_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06008_ _01512_ _01517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12605__CLK clknet_leaf_196_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11564__I0 _05713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09509__I0 _04371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08980__I1 u2.mem\[20\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07959_ u2.mem\[16\]\[15\] _03264_ _03265_ u2.mem\[33\]\[15\] _03423_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10119__I1 u2.mem\[46\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_2_0__f_clock_a_I clknet_0_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12755__CLK clknet_leaf_64_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10970_ _05360_ _01071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11867__I1 u2.mem\[191\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08709__S _03942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09629_ _04471_ u2.mem\[35\]\[3\] _04522_ _04526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11135__S _05462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12640_ _00519_ clknet_leaf_172_clock u2.mem\[32\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12571_ _00450_ clknet_leaf_182_clock u2.mem\[28\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07448__B2 u2.mem\[38\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11522_ _05706_ _01277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12135__CLK clknet_leaf_37_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11453_ _05661_ _01253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10773__I _05231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09996__I0 _04709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10404_ _03687_ _05009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11384_ _05619_ _01226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13123_ _01002_ clknet_leaf_21_clock u2.mem\[62\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_17_clock_I clknet_5_2_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10335_ _04963_ _00833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12285__CLK clknet_leaf_185_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06974__A3 _02424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13054_ _00933_ clknet_leaf_259_clock u2.mem\[58\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10266_ _04889_ u2.mem\[50\]\[1\] _04923_ _04925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13530__CLK clknet_leaf_317_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11555__I0 _05719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12005_ net24 clknet_2_3__leaf_clock_a mem_address_trans\[0\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08420__I0 _03685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10197_ _04878_ _00780_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09074__I _04181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07923__A2 _03385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08971__I1 u2.mem\[20\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11307__I0 _05552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08619__S _03880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07136__B1 _02614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12907_ _00786_ clknet_leaf_221_clock u2.mem\[49\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07687__A1 u2.mem\[8\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10948__I _04134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07687__B2 u2.mem\[4\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11045__S _05404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12838_ _00717_ clknet_leaf_63_clock u2.mem\[44\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12087__D net36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12769_ _00648_ clknet_leaf_154_clock u2.mem\[40\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06290_ u2.mem\[153\]\[2\] _01708_ _01710_ u2.mem\[160\]\[2\] _01795_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_334_clock clknet_5_6_0_clock clknet_leaf_334_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_72_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08354__S _03711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06111__A1 _01615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput20 data_in_a[7] net20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10683__I _05173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput31 mem_address_a[7] net31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06662__A2 _02012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13060__CLK clknet_leaf_27_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput42 row_select_a[5] net42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09987__I0 _04700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12628__CLK clknet_leaf_97_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11794__I0 _05876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_349_clock clknet_5_4_0_clock clknet_leaf_349_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09980_ _04694_ u2.mem\[43\]\[5\] _04745_ _04747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08931_ _04081_ _00311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12778__CLK clknet_leaf_130_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08862_ _03705_ _04039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10124__S _04835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08411__I0 _03668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06178__A1 u2.mem\[191\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06178__B2 u2.mem\[179\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08962__I1 u2.mem\[20\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07813_ u2.mem\[14\]\[12\] _03123_ _03124_ u2.mem\[12\]\[12\] _03280_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08793_ _03912_ u2.mem\[16\]\[3\] _03990_ _03994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07390__A3 _02853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07744_ u2.mem\[3\]\[11\] _03034_ _03211_ _03212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_42_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12008__CLK clknet_leaf_299_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07675_ _03141_ _03142_ _03143_ _03144_ _03145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10521__I1 u2.mem\[56\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09414_ _04393_ _04394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06626_ _02102_ _02106_ _02110_ _02111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09345_ _04272_ u2.mem\[28\]\[9\] _04346_ _04348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12158__CLK clknet_leaf_205_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08478__I0 _03719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06557_ _02041_ _02000_ _02042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09276_ _04281_ u2.mem\[26\]\[13\] _04305_ _04307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08264__S _03645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06102__A1 _01547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06488_ _01973_ _01970_ _01974_ _01975_ _01462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08227_ _03575_ u2.mem\[3\]\[13\] _03624_ _03626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06653__A2 _02136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09159__I _04225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09978__I0 _04691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08158_ _03539_ u2.mem\[2\]\[0\] _03585_ _03586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13553__CLK clknet_leaf_14_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11785__I0 _05870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07109_ u2.mem\[28\]\[0\] _02585_ _02587_ u2.mem\[31\]\[0\] _02588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08998__I _03987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08089_ data_in_trans\[15\].data_sync _03535_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09095__S _04192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10120_ _04833_ _00748_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06956__A3 _02433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10051_ _04788_ u2.mem\[45\]\[2\] _04784_ _04789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10034__S _04777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08012__B _03474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07407__I _02508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10969__S _05356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_243_clock_I clknet_5_19_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09622__I _04521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09902__I0 _04698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10953_ _05348_ _05349_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10512__I1 u2.mem\[56\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10884_ _05304_ _01041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12623_ _00502_ clknet_leaf_172_clock u2.mem\[31\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08469__I0 _03702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13083__CLK clknet_leaf_267_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12554_ _00433_ clknet_leaf_119_clock u2.mem\[26\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10976__A1 _04224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11505_ _05677_ u2.mem\[168\]\[4\] _05691_ _05697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12485_ _00364_ clknet_leaf_100_clock u2.mem\[22\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09969__I0 _04681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11436_ _05633_ u2.mem\[164\]\[4\] _05646_ _05652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08902__S _04061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11367_ _05587_ u2.mem\[160\]\[1\] _05608_ _05610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13106_ _00985_ clknet_leaf_241_clock u2.mem\[61\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10318_ _04943_ _04954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11298_ _05442_ _05566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13037_ _00916_ clknet_leaf_267_clock u2.mem\[57\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10249_ _04604_ _04913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07357__B1 _02674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07317__I _02456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06221__I _01726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07109__B1 _02587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08349__S _03711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11456__A2 _05645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12300__CLK clknet_leaf_181_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13426__CLK clknet_leaf_349_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07460_ u2.mem\[15\]\[6\] _02792_ _02793_ u2.mem\[13\]\[6\] _02933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06332__A1 u2.mem\[170\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07052__I _02530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06332__B2 u2.mem\[156\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06411_ u2.select_mem_row\[4\] u2.select_mem_col\[4\] _01502_ _01912_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07391_ _01843_ _02780_ _02820_ _02865_ _01496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_273_clock clknet_5_21_0_clock clknet_leaf_273_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_76_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11503__S _05692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09130_ _04154_ u2.mem\[23\]\[8\] _04213_ _04214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06342_ u2.mem\[189\]\[4\] _01650_ _01663_ u2.mem\[180\]\[4\] _01652_ u2.mem\[176\]\[4\]
+ _01845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__08085__A1 _01973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12450__CLK clknet_leaf_159_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13576__CLK clknet_leaf_32_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09061_ _04171_ u2.mem\[21\]\[13\] _04168_ _04172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10119__S _04830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06273_ _01625_ _01778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06635__A2 _02000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08880__I0 _04010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08012_ _01612_ _03471_ _03474_ _03475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_288_clock clknet_5_20_0_clock clknet_leaf_288_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_128_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_192_clock_I clknet_5_31_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11392__A1 _05295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06399__B2 u2.mem\[162\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_2_clock clknet_5_0_0_clock clknet_leaf_2_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09963_ _04714_ u2.mem\[42\]\[14\] _04734_ _04737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_211_clock clknet_5_29_0_clock clknet_leaf_211_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11519__I0 _05677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08914_ _04070_ _00305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09894_ _04693_ _00662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09643__S _04532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08845_ _04027_ _00279_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10789__S _05242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07899__B2 u2.mem\[21\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08776_ _03981_ _00256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_226_clock clknet_5_25_0_clock clknet_leaf_226_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_27_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06571__A1 u2.mem\[164\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06571__B2 u2.mem\[178\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input12_I data_in_a[14] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07727_ _03192_ _03193_ _03194_ _03195_ _03196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_2828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07658_ u2.mem\[49\]\[9\] _03126_ _03127_ u2.mem\[46\]\[9\] _03128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08058__I data_in_trans\[6\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06323__B2 u2.mem\[161\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07520__B1 _02900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06609_ _02093_ _02094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06874__A2 row_select_trans\[5\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07589_ u2.mem\[37\]\[8\] _03058_ _03059_ u2.mem\[59\]\[8\] _03060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11413__S _05638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09328_ _04338_ _00451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08076__A1 _03525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09259_ _04297_ _00423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10029__S _04772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12943__CLK clknet_leaf_237_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12270_ _00149_ clknet_leaf_185_clock u2.mem\[9\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08722__S _03947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11758__I0 _05835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11221_ _05354_ _05482_ _05519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_49_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11152_ _04071_ _05443_ _05474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_49_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10103_ _04790_ u2.mem\[46\]\[3\] _04820_ _04824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11083_ _05430_ u2.mem\[142\]\[4\] _05421_ _05431_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07339__B1 _02658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09553__S _04474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10034_ _04709_ u2.mem\[44\]\[12\] _04777_ _04778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10699__S _05184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11930__I0 _05211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11882__I _05928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12323__CLK clknet_leaf_84_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13449__CLK clknet_leaf_343_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06976__I _02454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10498__I _05050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11985_ _05990_ _01456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10936_ _04180_ _05317_ _05336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_90_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06314__A1 u2.mem\[172\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06314__B2 u2.mem\[180\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10867_ _05292_ _01036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11323__S _05575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12606_ _00485_ clknet_leaf_195_clock u2.mem\[30\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08067__A1 _03518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10798_ _05229_ u2.mem\[62\]\[15\] _05247_ _05251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_12537_ _00416_ clknet_leaf_116_clock u2.mem\[25\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07814__A1 u2.mem\[49\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06617__A2 _02100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07290__A2 _02580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12468_ _00347_ clknet_leaf_105_clock u2.mem\[21\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11419_ _05631_ u2.mem\[163\]\[3\] _05638_ _05642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12399_ _00278_ clknet_leaf_155_clock u2.mem\[17\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06960_ _02374_ _02439_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_136_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07047__I _02525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input4_I col_select_a[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06891_ _02369_ _02370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11921__I0 _05911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08630_ _03879_ _03890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07345__A3 _02812_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10402__S _05002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06553__A1 _02015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07896__A4 _03361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12816__CLK clknet_leaf_147_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06819__C _02299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08561_ _03824_ u2.mem\[10\]\[11\] _03846_ _03850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07512_ u2.mem\[58\]\[7\] _02809_ _02810_ u2.mem\[36\]\[7\] _02984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_139_clock_I clknet_5_13_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08492_ _03805_ _00148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08807__S _04000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07443_ u2.mem\[52\]\[5\] _02847_ _02848_ u2.mem\[21\]\[5\] _02917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_165_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06856__A2 _02329_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11233__S _05519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07374_ u2.mem\[52\]\[4\] _02847_ _02848_ u2.mem\[21\]\[4\] _02849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09113_ _04204_ _00370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06325_ u2.mem\[144\]\[3\] _01671_ _01673_ u2.mem\[182\]\[3\] _01829_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06608__A2 _02070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09044_ _04158_ u2.mem\[21\]\[9\] _04155_ _04159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09638__S _04527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06256_ u2.mem\[148\]\[1\] _01715_ _01698_ u2.mem\[154\]\[1\] u2.mem\[162\]\[1\]
+ _01700_ _01762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__06126__I _01632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11990__CLK clknet_leaf_329_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10871__I _03582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08605__I0 _03831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06187_ _01693_ _01694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_150_clock clknet_5_25_0_clock clknet_leaf_150_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_2_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10412__I0 _05014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08341__I _03708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07033__A2 _02509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12346__CLK clknet_leaf_59_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06241__B1 _01623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09946_ _04727_ _00680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06792__A1 u2.mem\[151\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06792__B2 u2.mem\[158\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_165_clock clknet_5_26_0_clock clknet_leaf_165_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_4016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09877_ _04564_ _04681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08828_ _04010_ u2.mem\[17\]\[0\] _04015_ _04016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10312__S _04949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06544__A1 _02023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12496__CLK clknet_leaf_163_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07741__B1 _03029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08759_ _03921_ u2.mem\[15\]\[7\] _03968_ _03972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11770_ _05833_ u2.mem\[185\]\[3\] _05857_ _05861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10721_ _04997_ _05202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06847__A2 _02128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13440_ _01319_ clknet_leaf_341_clock u2.mem\[176\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09097__I0 _04161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08516__I _03701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10652_ _05110_ u2.mem\[59\]\[7\] _05157_ _05161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_103_clock clknet_5_11_0_clock clknet_leaf_103_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_139_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07420__I _02532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13371_ _01250_ clknet_leaf_357_clock u2.mem\[165\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10982__S _05365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08844__I0 _04026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10583_ _05119_ u2.mem\[57\]\[11\] _05113_ _05120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12322_ _00201_ clknet_leaf_158_clock u2.mem\[12\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07272__A2 _02645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13121__CLK clknet_leaf_314_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11877__I _05928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12253_ _00132_ clknet_leaf_213_clock u2.mem\[8\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_118_clock clknet_5_15_0_clock clknet_leaf_118_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_141_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11204_ _05506_ _01159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12184_ _00063_ clknet_leaf_59_clock u2.mem\[3\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11135_ _05460_ u2.mem\[146\]\[0\] _05462_ _05463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13271__CLK clknet_leaf_5_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12839__CLK clknet_leaf_135_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11066_ _05392_ u2.mem\[141\]\[5\] _05412_ _05419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10017_ _04768_ _00710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_140_clock_I clknet_5_13_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12989__CLK clknet_leaf_258_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11968_ _05981_ _01448_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10095__A1 _04394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10956__I _04143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10919_ _05325_ _01055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11899_ _05941_ _01419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12219__CLK clknet_leaf_217_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06302__A4 _01806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09088__I0 _04148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13569_ _01448_ clknet_leaf_14_clock u2.mem\[194\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09458__S _04419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06110_ _01616_ _01617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07090_ _02566_ _02567_ _02425_ _02568_ _02569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_51_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11787__I _03670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12369__CLK clknet_leaf_223_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06041_ col_select_trans\[2\].data_sync col_select_trans\[3\].data_sync _01548_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11347__A1 _04417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09260__I0 _04265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_65_clock_I clknet_5_9_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09800_ _04615_ u2.mem\[38\]\[15\] _04633_ _04637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_82_clock clknet_5_9_0_clock clknet_leaf_82_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_87_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07992_ _03452_ _03453_ _03454_ _03455_ _03456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06774__A1 u2.mem\[168\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09193__S _04252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09731_ data_in_trans\[8\].data_sync _04591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06943_ _01551_ _02016_ _02422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09662_ _04545_ _00578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06874_ _01989_ row_select_trans\[5\].data_sync _02353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_95_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07723__B1 _03147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_97_clock clknet_5_10_0_clock clknet_leaf_97_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08613_ _03798_ u2.mem\[12\]\[0\] _03880_ _03881_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09593_ _04505_ _00549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08544_ _03840_ _00165_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09315__I1 u2.mem\[27\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08537__S _03836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09720__I _04582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11122__I1 u2.mem\[145\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08475_ _03794_ _00142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_20_clock clknet_5_2_0_clock clknet_leaf_20_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_165_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07426_ _02560_ _02900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09079__I0 _04132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13144__CLK clknet_leaf_39_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11898__S _05937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07357_ u2.mem\[26\]\[4\] _02673_ _02674_ u2.mem\[10\]\[4\] _02832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_342_clock_I clknet_5_5_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10633__I0 _05128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06308_ u2.mem\[171\]\[3\] _01611_ _01770_ u2.mem\[157\]\[3\] _01812_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_35_clock clknet_5_3_0_clock clknet_leaf_35_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_136_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07254__A2 _02687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07288_ u2.mem\[26\]\[3\] _02673_ _02674_ u2.mem\[10\]\[3\] _02764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09027_ _04145_ u2.mem\[21\]\[5\] _04141_ _04146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13294__CLK clknet_leaf_364_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06239_ _01738_ _01739_ _01744_ _01745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10307__S _04944_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11189__I1 u2.mem\[149\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09251__I0 _04256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06765__A1 u2.mem\[153\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07962__B1 _02505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06765__B2 u2.mem\[160\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09929_ _04717_ _00673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11138__S _05462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12940_ _00819_ clknet_leaf_256_clock u2.mem\[51\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07714__B1 _03056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09831__S _04654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12871_ _00750_ clknet_leaf_136_clock u2.mem\[46\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09306__I1 u2.mem\[27\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11822_ _05893_ _01390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08447__S _03778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11753_ _05851_ _01363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10704_ _05124_ u2.mem\[60\]\[13\] _05189_ _05191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11684_ _05768_ _05808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13423_ _01302_ clknet_leaf_348_clock u2.mem\[174\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10635_ _04311_ _05071_ _05151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__12511__CLK clknet_leaf_162_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11601__S _05747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09278__S _04305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10624__I0 _05119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13354_ _01233_ clknet_leaf_359_clock u2.mem\[162\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07245__A2 _02565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08182__S _03595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10566_ _03683_ _05108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12305_ _00184_ clknet_leaf_164_clock u2.mem\[11\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13285_ _01164_ clknet_leaf_0_clock u2.mem\[151\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10497_ _05065_ _00893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12236_ _00115_ clknet_leaf_211_clock u2.mem\[7\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12661__CLK clknet_leaf_77_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12167_ _00046_ clknet_leaf_109_clock u2.mem\[2\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06756__A1 _02209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11118_ _05285_ _05443_ _05452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_42_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12098_ _01496_ clknet_leaf_224_clock u2.active_mem\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13017__CLK clknet_leaf_319_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11049_ _05390_ u2.mem\[140\]\[4\] _05403_ _05409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 data_in_a[0] net7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07181__A1 u2.mem\[14\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_291_clock_I clknet_5_20_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12041__CLK clknet_2_3__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06590_ _02007_ _02037_ _02075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13167__CLK clknet_leaf_263_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08260_ _03566_ u2.mem\[4\]\[9\] _03645_ _03647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07211_ u2.mem\[5\]\[1\] _02687_ _02688_ u2.mem\[38\]\[1\] _02689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08191_ _03579_ u2.mem\[2\]\[15\] _03600_ _03604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12191__CLK clknet_leaf_237_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11511__S _05700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07142_ _02458_ _02459_ _02507_ _02364_ _02621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_9_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10615__I0 _05110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07236__A2 _02515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07073_ _02440_ _02378_ _02421_ _02552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_146_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06024_ u2.driver_mem\[8\] _01517_ _01532_ _01520_ _01533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_138_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07539__A3 _03009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07975_ u2.mem\[37\]\[15\] _03291_ _03292_ u2.mem\[59\]\[15\] _03439_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_45_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09714_ _04138_ _04578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06926_ _02398_ _02399_ _02400_ _02404_ _02405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_132_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09645_ _04487_ u2.mem\[35\]\[10\] _04532_ _04535_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06857_ _02309_ _02314_ _02323_ _02336_ _02337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_71_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09576_ _04494_ u2.mem\[33\]\[13\] _04492_ _04495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_06788_ _02266_ _02267_ _02268_ _02269_ _02270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_42_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08527_ _03829_ u2.mem\[9\]\[13\] _03827_ _03830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12534__CLK clknet_leaf_97_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08458_ _03681_ u2.mem\[8\]\[5\] _03783_ _03785_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08066__I _03493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07475__A2 _02937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07409_ u2.mem\[54\]\[5\] _02881_ _02882_ u2.mem\[55\]\[5\] _02883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08389_ _03706_ u2.mem\[6\]\[11\] _03738_ _03742_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11421__S _05637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10420_ _03708_ _05020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10606__I0 _05101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12684__CLK clknet_leaf_193_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10351_ _04973_ _00839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09826__S _04649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13070_ _00949_ clknet_leaf_253_clock u2.mem\[59\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10282_ _04904_ u2.mem\[50\]\[8\] _04933_ _04934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12021_ net32 clknet_2_1__leaf_clock_a mem_address_trans\[8\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06738__A1 u2.mem\[151\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07935__B1 _02575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06738__B2 u2.mem\[158\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09527__I1 u2.mem\[32\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07950__A3 _03409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12064__CLK clknet_leaf_300_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07145__I _02623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12923_ _00802_ clknet_leaf_252_clock u2.mem\[50\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12854_ _00733_ clknet_leaf_80_clock u2.mem\[45\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09360__I _04118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_13_clock_I clknet_5_3_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11098__I0 _05430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11805_ _05883_ _01383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12785_ _00664_ clknet_leaf_235_clock u2.mem\[41\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10845__I0 _05198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11736_ _05841_ _01356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07466__A2 _02881_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10470__A1 _03752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11667_ _05679_ _05798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_168_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13406_ _01285_ clknet_leaf_304_clock u2.mem\[171\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07218__A2 _02633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10618_ _05112_ u2.mem\[58\]\[8\] _05141_ _05142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11598_ _05754_ u2.mem\[174\]\[3\] _05748_ _05755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11270__I0 _05548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_238_clock_I clknet_5_19_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13337_ _01216_ clknet_leaf_9_clock u2.mem\[159\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10549_ _05096_ _00914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06977__A1 _02451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09215__I0 _04267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13268_ _01147_ clknet_leaf_9_clock u2.mem\[148\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11022__I0 _05392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12219_ _00098_ clknet_leaf_217_clock u2.mem\[6\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13199_ _01078_ clknet_leaf_274_clock u2.mem\[136\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06729__A1 u2.mem\[176\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07926__B1 _02533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06729__B2 u2.mem\[189\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12407__CLK clknet_leaf_112_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09518__I1 u2.mem\[32\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07760_ u2.mem\[57\]\[11\] _03061_ _03062_ u2.mem\[41\]\[11\] _03228_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06711_ u2.mem\[154\]\[1\] _02126_ _02129_ u2.mem\[148\]\[1\] _02127_ u2.mem\[162\]\[1\]
+ _02195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_38_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07691_ _01958_ _03013_ _03131_ _03160_ _01501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07154__A1 _01544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12557__CLK clknet_leaf_192_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09430_ _04371_ u2.mem\[30\]\[6\] _04401_ _04404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06642_ _02007_ _02052_ _02127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06901__A1 _02352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09361_ _03904_ _04250_ _04357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06573_ _02026_ _02036_ _02058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08312_ _03685_ u2.mem\[5\]\[6\] _03677_ _03686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09292_ _04258_ u2.mem\[27\]\[3\] _04313_ _04317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08243_ _03637_ _00067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08174_ _03594_ _00041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07125_ u2.mem\[52\]\[0\] _02601_ _02603_ u2.mem\[21\]\[0\] _02604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06968__A1 _02429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11040__I _05403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07056_ _02518_ _02524_ _02529_ _02534_ _02535_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09206__I0 _04260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11975__I _05970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11013__I0 _05386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06007_ u2.select_mem_row\[2\] u2.select_mem_col\[2\] _01510_ _01516_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12087__CLK clknet_2_1__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input42_I row_select_a[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09509__I1 u2.mem\[32\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07958_ u2.mem\[1\]\[15\] _03261_ _03262_ u2.mem\[7\]\[15\] _03422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06909_ _02387_ _02388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_99_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07889_ u2.mem\[37\]\[13\] _03291_ _03292_ u2.mem\[59\]\[13\] _03355_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13482__CLK clknet_leaf_298_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09628_ _04525_ _00564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_187_clock_I clknet_5_31_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09559_ _04464_ _04483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_24_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12570_ _00449_ clknet_leaf_111_clock u2.mem\[27\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07448__A2 _02920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11521_ _05680_ u2.mem\[169\]\[5\] _05699_ _05706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11452_ _05635_ u2.mem\[165\]\[5\] _05654_ _05661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10403_ _05008_ _00856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11383_ _05589_ u2.mem\[161\]\[2\] _05616_ _05619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09556__S _04474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06044__I col_select_trans\[4\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13122_ _01001_ clknet_leaf_242_clock u2.mem\[62\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10334_ _04920_ u2.mem\[51\]\[15\] _04959_ _04963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08460__S _03783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13053_ _00932_ clknet_leaf_259_clock u2.mem\[58\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06979__I _02417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10265_ _04924_ _00802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11555__I1 u2.mem\[171\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12004_ _00016_ clknet_leaf_40_clock u2.mem\[0\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10196_ _04806_ u2.mem\[48\]\[10\] _04875_ _04878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11307__I1 u2.mem\[156\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12906_ _00785_ clknet_leaf_141_clock u2.mem\[48\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07687__A2 _03091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12837_ _00716_ clknet_leaf_82_clock u2.mem\[44\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12768_ _00647_ clknet_leaf_155_clock u2.mem\[40\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08635__S _03890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11719_ _05829_ u2.mem\[182\]\[1\] _05827_ _05830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13205__CLK clknet_leaf_275_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12699_ _00578_ clknet_leaf_255_clock u2.mem\[36\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06111__A2 _01617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput10 data_in_a[12] net10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 data_in_a[8] net21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput32 mem_address_a[8] net32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05994__S _01502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11794__I1 u2.mem\[186\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07611__A2 _03080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13355__CLK clknet_leaf_360_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08930_ _04026_ u2.mem\[19\]\[5\] _04079_ _04081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06889__I _02353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10405__S _05002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08861_ _04038_ _00284_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07812_ u2.mem\[44\]\[12\] _03120_ _03121_ u2.mem\[42\]\[12\] _03279_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08792_ _03993_ _00260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07743_ _02357_ _03211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07390__A4 _02864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07674_ u2.mem\[28\]\[9\] _03072_ _03073_ u2.mem\[31\]\[9\] _03144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10140__S _04841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07678__A2 _03146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06625_ u2.mem\[159\]\[0\] _02107_ _02109_ u2.mem\[149\]\[0\] _02110_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09413_ _03581_ _03902_ _04393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_164_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06350__A2 _01850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09344_ _04347_ _00458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06556_ _02036_ _02001_ _02041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06129__I _01635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09275_ _04306_ _00430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11482__I0 _05663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06487_ u2.mem\[193\]\[13\] _01917_ _01919_ u2.mem\[192\]\[13\] _01964_ _01975_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_32_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08226_ _03625_ _00062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08157_ _03584_ _03585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_107_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07108_ _02586_ _02587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08088_ _01976_ _03527_ _03534_ _00015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07039_ u2.mem\[43\]\[0\] _02515_ _02517_ u2.mem\[20\]\[0\] _02518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06956__A4 _02434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12722__CLK clknet_leaf_235_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10050_ _04572_ _04788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07366__A1 u2.mem\[28\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10114__I _04819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08519__I _03705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10952_ _04138_ _05348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10673__A1 _04334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13228__CLK clknet_leaf_280_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10883_ _05303_ u2.mem\[130\]\[3\] _05297_ _05304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12622_ _00501_ clknet_leaf_189_clock u2.mem\[31\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12553_ _00432_ clknet_leaf_119_clock u2.mem\[26\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11504_ _05696_ _01269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12252__CLK clknet_leaf_215_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12484_ _00363_ clknet_leaf_105_clock u2.mem\[22\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13378__CLK clknet_leaf_36_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11435_ _05651_ _01245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09286__S _04313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11366_ _05609_ _01218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10317_ _04953_ _00825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13105_ _00984_ clknet_leaf_314_clock u2.mem\[61\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10225__S _04896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11297_ _05565_ _01193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10248_ _04912_ _00797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13036_ _00915_ clknet_leaf_260_clock u2.mem\[57\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07357__B2 u2.mem\[10\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10024__I _04761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10179_ _04868_ _00772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07109__B2 u2.mem\[31\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11056__S _05413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06580__A2 _02028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10895__S _05310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06410_ u2.select_mem_row\[5\] u2.select_mem_col\[5\] _01510_ _01911_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07390_ _02831_ _02842_ _02853_ _02864_ _02865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_22_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08365__S _03728_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06341_ _01843_ _01844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06096__A1 _01566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09060_ _04170_ _04171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07293__B1 _02681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06272_ u2.mem\[167\]\[2\] _01775_ _01776_ u2.mem\[183\]\[2\] _01777_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08011_ _03472_ _03473_ _01549_ _03474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12745__CLK clknet_leaf_53_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09196__S _04252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07045__B1 _02523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_135_clock_I clknet_5_13_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06399__A2 _01699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11392__A2 _05606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09962_ _04736_ _00687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11519__I1 u2.mem\[169\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08913_ _04048_ u2.mem\[18\]\[15\] _04066_ _04070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09893_ _04691_ u2.mem\[41\]\[4\] _04692_ _04693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08396__I0 _03719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08844_ _04026_ u2.mem\[17\]\[5\] _04024_ _04027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09723__I data_in_trans\[6\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06020__A1 u2.driver_mem\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08775_ _03937_ u2.mem\[15\]\[14\] _03978_ _03981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08148__I0 _03577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07726_ u2.mem\[18\]\[10\] _03083_ _03084_ u2.mem\[19\]\[10\] _03195_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09896__I0 _04694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07657_ _02532_ _03127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06608_ _02031_ _02070_ _02093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12275__CLK clknet_leaf_102_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07588_ _02541_ _03059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13520__CLK clknet_leaf_16_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09327_ _04254_ u2.mem\[28\]\[1\] _04336_ _04338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06539_ row_select_trans\[1\].data_sync _02024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_139_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08076__A2 _03519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06087__A1 _01556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07284__B1 _02549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09258_ _04263_ u2.mem\[26\]\[5\] _04295_ _04297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08209_ _03557_ u2.mem\[3\]\[5\] _03614_ _03616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09189_ _04248_ _04249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_135_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11220_ _05518_ _01163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11758__I1 u2.mem\[184\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11151_ _05473_ _01139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10045__S _04784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07051__A3 _02433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10102_ _04823_ _00740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11082_ _05348_ _05430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07339__B2 u2.mem\[12\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08387__I0 _03702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10033_ _04761_ _04777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_114_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08000__A2 _03461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10194__I0 _04804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_333_clock clknet_5_6_0_clock clknet_leaf_333_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_76_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_337_clock_I clknet_5_4_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13050__CLK clknet_leaf_44_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11984_ _05227_ u2.mem\[194\]\[14\] _05971_ _05990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12618__CLK clknet_leaf_111_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10935_ _05334_ _05335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_348_clock clknet_5_4_0_clock clknet_leaf_348_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_147_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06314__A2 _01654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11604__S _05747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06992__I _02470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08185__S _03600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10866_ _05204_ u2.mem\[129\]\[4\] _05286_ _05292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12605_ _00484_ clknet_leaf_196_clock u2.mem\[30\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11446__I0 _05629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08067__A2 _03519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12768__CLK clknet_leaf_155_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10797_ _05250_ _01008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_12536_ _00415_ clknet_leaf_116_clock u2.mem\[25\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07102__B _02552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08913__S _04066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07814__A2 _03126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12467_ _00346_ clknet_leaf_108_clock u2.mem\[21\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07027__B1 _02505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11418_ _05641_ _01238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12398_ _00277_ clknet_leaf_179_clock u2.mem\[17\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11349_ _05583_ u2.mem\[159\]\[0\] _05598_ _05599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06786__C1 u2.mem\[144\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06250__A1 u2.mem\[187\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06250__B2 u2.mem\[192\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12148__CLK clknet_leaf_74_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08378__I0 _03685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13019_ _00898_ clknet_leaf_249_clock u2.mem\[56\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06890_ _02366_ _02367_ _02368_ _02369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_45_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10185__I0 _04795_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11921__I1 u2.mem\[193\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07345__A4 _02819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06553__A2 _02037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08560_ _03849_ _00172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12298__CLK clknet_leaf_165_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07063__I _02541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13543__CLK clknet_leaf_32_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07511_ u2.mem\[53\]\[7\] _02806_ _02807_ u2.mem\[56\]\[7\] _02983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08491_ _03804_ u2.mem\[9\]\[2\] _03800_ _03805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08550__I0 _03813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07998__I _01547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07442_ u2.mem\[17\]\[5\] _02844_ _02845_ u2.mem\[24\]\[5\] _02916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_61_clock_I clknet_5_9_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07373_ _02602_ _02848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08302__I0 _03676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09112_ _04119_ u2.mem\[23\]\[0\] _04203_ _04204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06324_ _01820_ _01821_ _01822_ _01827_ _01828_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07266__B1 _02461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09043_ _04157_ _04158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06255_ u2.mem\[152\]\[1\] _01713_ _01708_ u2.mem\[153\]\[1\] _01761_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_11_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06186_ _01563_ _01677_ _01580_ _01693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA_clkbuf_leaf_286_clock_I clknet_5_20_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_13_0_clock clknet_3_6_0_clock clknet_4_13_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_150_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06241__A1 u2.mem\[167\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09945_ _04696_ u2.mem\[42\]\[6\] _04724_ _04727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06241__B2 u2.mem\[183\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08369__I0 _03668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06792__A2 _02084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13073__CLK clknet_leaf_236_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09876_ _04680_ _00657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10176__I0 _04786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09453__I _04416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08827_ _04014_ _04015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_3305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10599__I _05130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06544__A2 _02028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08069__I data_in_trans\[9\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08758_ _03971_ _00248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09869__I0 _04605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07709_ u2.mem\[49\]\[10\] _03126_ _03127_ u2.mem\[46\]\[10\] _03178_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11676__I0 _05792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09494__A1 _03983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08689_ _03705_ _03930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08541__I0 _03804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12910__CLK clknet_leaf_202_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10720_ _05201_ _00980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11428__I0 _05623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10651_ _05160_ _00952_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07257__B1 _02624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13370_ _01249_ clknet_leaf_357_clock u2.mem\[165\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10582_ _03704_ _05119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12321_ _00200_ clknet_leaf_158_clock u2.mem\[12\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10800__A1 _04416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08532__I _03722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12252_ _00131_ clknet_leaf_215_clock u2.mem\[8\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11203_ _05505_ u2.mem\[150\]\[1\] _05502_ _05506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12183_ _00062_ clknet_leaf_61_clock u2.mem\[3\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13416__CLK clknet_leaf_341_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07148__I _02626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06232__A1 u2.mem\[144\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06232__B2 u2.mem\[182\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06052__I col_select_trans\[3\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11134_ _05461_ _05462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07980__A1 u2.mem\[9\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_272_clock clknet_5_20_0_clock clknet_leaf_272_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_95_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07980__B2 u2.mem\[25\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11065_ _05418_ _01108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10167__I0 _04817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06987__I _02387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10503__S _05066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12440__CLK clknet_leaf_123_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10016_ _04691_ u2.mem\[44\]\[4\] _04767_ _04768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11903__I1 _03525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13566__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_287_clock clknet_5_20_0_clock clknet_leaf_287_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11967_ _05209_ u2.mem\[194\]\[6\] _05980_ _05981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12590__CLK clknet_leaf_190_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10095__A2 _04760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_1_clock clknet_5_0_0_clock clknet_leaf_1_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10918_ _05307_ u2.mem\[132\]\[5\] _05318_ _05325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11898_ u2.mem\[192\]\[9\] _03521_ _05937_ _05941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_210_clock clknet_5_29_0_clock clknet_leaf_210_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11419__I0 _05631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10849_ _05202_ u2.mem\[128\]\[3\] _05278_ _05282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13568_ _01447_ clknet_leaf_15_clock u2.mem\[194\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12519_ _00398_ clknet_leaf_117_clock u2.mem\[24\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13499_ _01378_ clknet_leaf_316_clock u2.mem\[186\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_225_clock clknet_5_25_0_clock clknet_leaf_225_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_12_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06040_ _01546_ _01547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07058__I _02370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_21_0_clock_I clknet_4_10_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07991_ u2.mem\[6\]\[15\] _03327_ _03328_ u2.mem\[47\]\[15\] _03455_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06774__A2 _02093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09730_ _04590_ _00601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10158__I0 _04808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06942_ _02402_ _02421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_79_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09273__I _04289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09661_ _04463_ u2.mem\[36\]\[0\] _04544_ _04545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06873_ _02340_ _02352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08771__I0 _03932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08612_ _03879_ _03880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_23_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12933__CLK clknet_leaf_67_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09592_ _04471_ u2.mem\[34\]\[3\] _04501_ _04505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08543_ _03806_ u2.mem\[10\]\[3\] _03836_ _03840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08279__A2 _03544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11244__S _05529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08474_ _03710_ u2.mem\[8\]\[12\] _03793_ _03794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10330__I0 _04916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06829__A3 _02307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07425_ _02558_ _02899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07239__B1 _02667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07356_ _02821_ _02824_ _02827_ _02830_ _02831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_149_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06307_ u2.mem\[167\]\[3\] _01775_ _01776_ u2.mem\[183\]\[3\] _01811_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10882__I _04997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12313__CLK clknet_leaf_118_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07287_ _02759_ _02760_ _02761_ _02762_ _02763_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__13439__CLK clknet_leaf_341_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09026_ _04144_ _04145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06238_ u2.mem\[147\]\[1\] _01676_ _01680_ u2.mem\[169\]\[1\] _01743_ _01744_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_156_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08352__I _03717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06169_ _01675_ _01676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09251__I1 u2.mem\[26\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06214__A1 _01678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12463__CLK clknet_leaf_172_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11419__S _05638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10323__S _04954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09928_ _04716_ u2.mem\[41\]\[15\] _04710_ _04717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10149__I0 _04799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06600__I _02084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09859_ _04660_ _04671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_115_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08762__I0 _03923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11218__I _05516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12870_ _00749_ clknet_leaf_83_clock u2.mem\[46\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07190__A2 _02666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11821_ _05874_ u2.mem\[188\]\[4\] _05887_ _05893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08514__I0 _03820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11752_ _05829_ u2.mem\[184\]\[1\] _05849_ _05851_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10321__I0 _04907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10703_ _05190_ _00974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11683_ _05807_ _01337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13422_ _01301_ clknet_leaf_309_clock u2.mem\[173\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06047__I _01553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10634_ _05150_ _00945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13353_ _01232_ clknet_leaf_358_clock u2.mem\[162\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11821__I0 _05874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10565_ _05107_ _00919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12304_ _00183_ clknet_leaf_164_clock u2.mem\[11\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13284_ _01163_ clknet_leaf_1_clock u2.mem\[150\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10496_ _05018_ u2.mem\[55\]\[11\] _05061_ _05065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12235_ _00114_ clknet_leaf_211_clock u2.mem\[7\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12166_ _00045_ clknet_leaf_91_clock u2.mem\[2\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06756__A2 _02214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11117_ _05451_ _01127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12956__CLK clknet_leaf_197_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12097_ _01495_ clknet_leaf_219_clock u2.active_mem\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07606__I _02590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11048_ _05408_ _01101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07705__A1 u2.mem\[58\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput8 data_in_a[10] net8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08753__I0 _03914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07705__B2 u2.mem\[36\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_234_clock_I clknet_5_18_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07181__A2 _02657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09821__I _04638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12999_ _00878_ clknet_leaf_323_clock u2.mem\[54\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11064__S _05412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11265__A1 _04287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10312__I0 _04898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07341__I _02514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07210_ _02628_ _02688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08190_ _03603_ _00048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_164_clock clknet_5_26_0_clock clknet_leaf_164_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07141_ u2.mem\[39\]\[0\] _02617_ _02619_ u2.mem\[48\]\[0\] _02620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10615__I1 u2.mem\[58\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06444__A1 _01844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12486__CLK clknet_leaf_100_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07072_ _02347_ _02551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_145_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06023_ u2.driver_mem\[9\] _01518_ _01532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_86_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_179_clock clknet_5_30_0_clock clknet_leaf_179_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_160_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07944__A1 _03405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07974_ u2.mem\[60\]\[15\] _03288_ _03289_ u2.mem\[62\]\[15\] _03438_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_19_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_102_clock clknet_5_11_0_clock clknet_leaf_102_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09932__S _04719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09713_ _04577_ _00597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06925_ _02401_ _02403_ _02383_ _02404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_19_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08744__I0 _03900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11038__I _05275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09644_ _04534_ _00571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07960__B _02358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06856_ _02324_ _02329_ _02330_ _02335_ _02336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_56_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10551__I0 _05097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09731__I data_in_trans\[8\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13111__CLK clknet_leaf_38_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07172__A2 _02648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09575_ _04170_ _04494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_06787_ u2.mem\[146\]\[3\] _02156_ _02122_ u2.mem\[173\]\[3\] _02269_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_117_clock clknet_5_14_0_clock clknet_leaf_117_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_97_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08526_ _03714_ _03829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10303__I0 _04889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08347__I _03713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08457_ _03784_ _00134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07475__A3 _02942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13261__CLK clknet_leaf_270_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06683__A1 u2.mem\[170\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07408_ _02510_ _02882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06683__B2 u2.mem\[156\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08388_ _03741_ _00108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12829__CLK clknet_leaf_207_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07339_ u2.mem\[14\]\[4\] _02657_ _02658_ u2.mem\[12\]\[4\] _02814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09621__A1 _04072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10350_ _04898_ u2.mem\[52\]\[5\] _04971_ _04973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09009_ _04130_ _04131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10281_ _04922_ _04933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_69_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12979__CLK clknet_leaf_42_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_183_clock_I clknet_5_30_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12020_ mem_address_trans\[7\].A clknet_leaf_289_clock mem_address_trans\[7\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06199__B1 _01705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07935__B2 u2.mem\[10\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12209__CLK clknet_leaf_232_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07426__I _02560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09842__S _04661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10988__S _05364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07950__A4 _03414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12922_ _00801_ clknet_leaf_126_clock u2.mem\[49\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11495__A1 _04223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07699__B1 _03032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08458__S _03783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12853_ _00732_ clknet_leaf_80_clock u2.mem\[45\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12359__CLK clknet_leaf_133_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06371__B1 _01679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11804_ _05872_ u2.mem\[187\]\[3\] _05879_ _05883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08257__I _03634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12784_ _00663_ clknet_leaf_321_clock u2.mem\[41\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09160__I0 _04140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11735_ _05825_ u2.mem\[183\]\[0\] _05840_ _05841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_81_clock clknet_5_8_0_clock clknet_leaf_81_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_41_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11612__S _05761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06674__A1 u2.mem\[146\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06674__B2 u2.mem\[186\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10470__A2 _04964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11666_ _05797_ _01330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13405_ _01284_ clknet_leaf_304_clock u2.mem\[171\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10617_ _05130_ _05141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10228__S _04896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11597_ _05673_ _05754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_155_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06426__A1 u2.mem\[194\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13336_ _01215_ clknet_leaf_17_clock u2.mem\[159\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_96_clock clknet_5_10_0_clock clknet_leaf_96_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08921__S _04074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11270__I1 u2.mem\[154\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10548_ _05093_ u2.mem\[57\]\[0\] _05095_ _05096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06977__A2 _02452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13267_ _01146_ clknet_leaf_5_clock u2.mem\[148\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10479_ _05055_ _00885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12218_ _00097_ clknet_leaf_52_clock u2.mem\[5\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13198_ _01077_ clknet_leaf_276_clock u2.mem\[136\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07926__A1 u2.mem\[49\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12149_ _00028_ clknet_leaf_73_clock u2.mem\[1\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13134__CLK clknet_leaf_268_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06710_ _02191_ _02193_ _02194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07690_ _03138_ _03145_ _03152_ _03159_ _03160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_38_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_34_clock clknet_5_3_0_clock clknet_leaf_34_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07154__A2 _02361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06641_ _02045_ _02125_ _02126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_64_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06362__B1 _01715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09360_ _04118_ _04356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06572_ _02006_ _02057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09151__I0 _04119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08311_ _03684_ _03685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09291_ _04316_ _00436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_49_clock clknet_5_7_0_clock clknet_leaf_49_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_33_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09199__S _04252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08242_ _03548_ u2.mem\[4\]\[1\] _03635_ _03637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08173_ _03561_ u2.mem\[2\]\[7\] _03590_ _03594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10138__S _04841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06417__A1 _01911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07124_ _02602_ _02603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07614__B1 _03084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08831__S _04015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06415__I _01912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06968__A2 _02445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07055_ u2.mem\[49\]\[0\] _02531_ _02533_ u2.mem\[46\]\[0\] _02534_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09206__I1 u2.mem\[25\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06006_ _01504_ _01509_ _01514_ _01515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08630__I _03879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06150__I _01656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input35_I output_active_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07957_ u2.mem\[15\]\[15\] _03258_ _03259_ u2.mem\[13\]\[15\] _03421_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12501__CLK clknet_leaf_106_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06908_ _02365_ _02372_ _02353_ _02387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_83_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07888_ u2.mem\[60\]\[13\] _03288_ _03289_ u2.mem\[62\]\[13\] _03354_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_16_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09627_ _04469_ u2.mem\[35\]\[2\] _04522_ _04525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06839_ u2.mem\[166\]\[5\] _02097_ _02099_ u2.mem\[161\]\[5\] _02318_ _02319_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_55_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06353__B1 _01734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09558_ _04153_ _04482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_169_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12651__CLK clknet_leaf_207_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08509_ _03692_ _03817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09489_ _04391_ u2.mem\[31\]\[15\] _04434_ _04438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11520_ _05705_ _01276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07853__B1 _03154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11451_ _05660_ _01252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13007__CLK clknet_leaf_240_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10048__S _04784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06408__A1 _01882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09837__S _04654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10402_ _05007_ u2.mem\[53\]\[6\] _05002_ _05008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07605__B1 _02914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11252__I1 u2.mem\[153\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11382_ _05618_ _01225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07081__A1 _02473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13121_ _01000_ clknet_leaf_314_clock u2.mem\[62\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10333_ _04962_ _00832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12031__CLK clknet_2_3__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13052_ _00931_ clknet_leaf_259_clock u2.mem\[58\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10264_ _04885_ u2.mem\[50\]\[0\] _04923_ _04924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07908__A1 _01973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12003_ _00015_ clknet_leaf_41_clock u2.mem\[0\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10195_ _04877_ _00779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07156__I _02447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06060__I _01566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12181__CLK clknet_leaf_77_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09371__I _04135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07136__A2 _02612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12905_ _00784_ clknet_leaf_141_clock u2.mem\[48\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12836_ _00715_ clknet_leaf_61_clock u2.mem\[44\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07105__B _02519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12767_ _00646_ clknet_leaf_155_clock u2.mem\[40\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11342__S _05584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06647__A1 u2.mem\[148\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06647__B2 u2.mem\[152\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11718_ _03662_ _05829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08715__I _03941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12698_ _00577_ clknet_leaf_110_clock u2.mem\[35\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput11 data_in_a[13] net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11649_ _05785_ _01325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput22 data_in_a[9] net22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput33 mem_address_a[9] net33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13319_ _01198_ clknet_leaf_301_clock u2.mem\[156\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09546__I _04464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12524__CLK clknet_leaf_187_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08860_ _04037_ u2.mem\[17\]\[10\] _04033_ _04038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08572__A1 _03605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07811_ _03270_ _03271_ _03274_ _03277_ _03278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_57_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08791_ _03910_ u2.mem\[16\]\[2\] _03990_ _03993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11517__S _05700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07742_ u2.mem\[16\]\[11\] _03031_ _03032_ u2.mem\[33\]\[11\] _03210_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09372__I0 _04364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12674__CLK clknet_leaf_154_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07673_ u2.mem\[9\]\[9\] _03069_ _03070_ u2.mem\[25\]\[9\] _03143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_4_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09412_ _04392_ _00481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_131_clock_I clknet_5_12_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06624_ _02108_ _02037_ _02109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09343_ _04269_ u2.mem\[28\]\[8\] _04346_ _04347_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06555_ u2.mem\[155\]\[0\] _02030_ _02035_ u2.mem\[174\]\[0\] u2.mem\[181\]\[0\]
+ _02039_ _02040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_33_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11252__S _05537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09274_ _04278_ u2.mem\[26\]\[12\] _04305_ _04306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11482__I1 u2.mem\[167\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06486_ u2.mem\[194\]\[13\] _01933_ _01974_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08225_ _03572_ u2.mem\[3\]\[12\] _03624_ _03625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12054__CLK clknet_leaf_287_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08561__S _03846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08156_ _03480_ _03583_ _03584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_162_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07107_ _02388_ _02390_ _02453_ _02473_ _02586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_101_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08087_ _03533_ _03529_ _03534_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06810__A1 u2.mem\[146\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07038_ _02516_ _02517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06810__B2 u2.mem\[186\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_56_clock_I clknet_5_12_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10745__I0 _05218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09392__S _04376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08989_ _04046_ u2.mem\[20\]\[14\] _04112_ _04115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09363__I0 _04356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06748__C _02230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10951_ _05347_ _01065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06326__B1 _01704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06877__A1 _02352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10882_ _04997_ _05303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12621_ _00500_ clknet_leaf_190_clock u2.mem\[31\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11162__S _05474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12552_ _00431_ clknet_leaf_119_clock u2.mem\[26\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11622__A1 _03487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06483__C _01964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11503_ _05674_ u2.mem\[168\]\[3\] _05692_ _05696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12483_ _00362_ clknet_leaf_123_clock u2.mem\[22\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_333_clock_I clknet_5_6_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11225__I1 u2.mem\[151\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11434_ _05631_ u2.mem\[164\]\[3\] _05647_ _05651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06055__I col_select_trans\[0\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08471__S _03788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12547__CLK clknet_leaf_103_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11365_ _05583_ u2.mem\[160\]\[0\] _05608_ _05609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10984__I0 _05346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13104_ _00983_ clknet_leaf_243_clock u2.mem\[61\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10316_ _04902_ u2.mem\[51\]\[7\] _04949_ _04953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06801__A1 u2.mem\[171\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06801__B2 u2.mem\[157\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11296_ _05556_ u2.mem\[155\]\[5\] _05558_ _05565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08003__B1 _03459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13035_ _00914_ clknet_leaf_248_clock u2.mem\[57\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10247_ _04911_ u2.mem\[49\]\[11\] _04905_ _04912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07357__A2 _02673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12697__CLK clknet_leaf_111_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10178_ _04788_ u2.mem\[48\]\[2\] _04865_ _04868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10241__S _04905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07109__A2 _02585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09354__I0 _04281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06317__C2 u2.mem\[193\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09106__I0 _04174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12819_ _00698_ clknet_leaf_60_clock u2.mem\[43\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10975__I _05275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12077__CLK clknet_2_2__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06340_ u2.mem\[0\]\[4\] _01843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_33_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13322__CLK clknet_leaf_342_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06393__C _01894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06271_ _01623_ _01776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06096__A2 _01599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08010_ u2.active_mem\[0\] _03458_ _03459_ u2.active_mem\[1\] _03473_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__11800__S _05879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06253__C1 _01660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09961_ _04712_ u2.mem\[42\]\[13\] _04734_ _04736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07060__A4 _02484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08912_ _04069_ _00304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09892_ _04682_ _04692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08843_ _03680_ _04026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08774_ _03980_ _00255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08148__I1 u2.mem\[1\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09345__I0 _04272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07725_ u2.mem\[52\]\[10\] _03080_ _03081_ u2.mem\[21\]\[10\] _03194_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_282_clock_I clknet_5_21_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07656_ _02530_ _03126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07520__A2 _02899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06607_ _02091_ _02092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10885__I _05000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07587_ _02539_ _03058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09326_ _04337_ _00450_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06538_ _02022_ _02023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09257_ _04296_ _00422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06469_ u2.mem\[193\]\[9\] _01960_ _01943_ u2.mem\[194\]\[9\] _01949_ _01961_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_166_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08208_ _03615_ _00054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08291__S _03660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11207__I1 u2.mem\[150\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09188_ _03901_ _04247_ _04248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_120_1566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08139_ _03571_ _00029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09186__I _04118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11150_ _05472_ u2.mem\[146\]\[5\] _05461_ _05473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07051__A4 _02463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10101_ _04788_ u2.mem\[46\]\[2\] _04820_ _04823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11081_ _05429_ _01113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07339__A2 _02657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10032_ _04776_ _00717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09336__I0 _04263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06478__C _01964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10996__S _05373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11983_ _05989_ _01455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10934_ _04117_ _05334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13345__CLK clknet_leaf_4_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10865_ _05291_ _01035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12604_ _00483_ clknet_leaf_191_clock u2.mem\[30\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11446__I1 u2.mem\[165\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_10796_ _05227_ u2.mem\[62\]\[14\] _05247_ _05250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12535_ _00414_ clknet_leaf_115_clock u2.mem\[25\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07102__C _02426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12466_ _00345_ clknet_leaf_162_clock u2.mem\[21\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11417_ _05629_ u2.mem\[163\]\[2\] _05638_ _05641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12397_ _00276_ clknet_leaf_180_clock u2.mem\[17\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07609__I _02600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11348_ _05597_ _05598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_98_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06786__B1 _02116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06786__C2 _02114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11279_ _05554_ u2.mem\[154\]\[4\] _05545_ _05555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13018_ _00897_ clknet_leaf_322_clock u2.mem\[55\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10185__I1 u2.mem\[48\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06002__A2 _01502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09327__I0 _04254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07510_ u2.mem\[54\]\[7\] _02881_ _02882_ u2.mem\[55\]\[7\] _02982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08490_ _03667_ _03804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08376__S _03733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08550__I1 u2.mem\[10\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07441_ u2.mem\[23\]\[5\] _02913_ _02914_ u2.mem\[22\]\[5\] _02915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12712__CLK clknet_leaf_50_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07372_ _02600_ _02847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08175__I _03584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09111_ _04202_ _04203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_149_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06323_ u2.mem\[166\]\[3\] _01753_ _01754_ u2.mem\[161\]\[3\] _01826_ _01827_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_104_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09042_ data_in_trans\[9\].data_sync _04157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06254_ u2.mem\[180\]\[1\] _01664_ _01666_ u2.mem\[150\]\[1\] _01760_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_15_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12862__CLK clknet_leaf_199_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_229_clock_I clknet_5_25_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06185_ _01691_ _01692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06423__I _01923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06777__B1 _02091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09944_ _04726_ _00679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13218__CLK clknet_leaf_283_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06241__A2 _01622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09566__I0 _04487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09875_ _04615_ u2.mem\[40\]\[15\] _04676_ _04680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11373__I0 _05593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09191__A1 _04249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08826_ _04011_ _04013_ _04014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12242__CLK clknet_leaf_226_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07741__A2 _03028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09670__S _04549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13368__CLK clknet_leaf_359_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08757_ _03919_ u2.mem\[15\]\[6\] _03968_ _03971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_1494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07708_ u2.mem\[14\]\[10\] _03123_ _03124_ u2.mem\[12\]\[10\] _03177_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11825__A1 _05411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08688_ _03929_ _00220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08286__S _03660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11676__I1 u2.mem\[179\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09494__A2 _04441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07639_ u2.mem\[3\]\[9\] _03034_ _02978_ _03109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12392__CLK clknet_leaf_133_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11428__I1 u2.mem\[164\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10650_ _05108_ u2.mem\[59\]\[6\] _05157_ _05160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09309_ _04326_ _00444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10581_ _05118_ _00924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12320_ _00199_ clknet_leaf_158_clock u2.mem\[12\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08813__I _03989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07009__A1 _02487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12251_ _00130_ clknet_leaf_216_clock u2.mem\[8\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11202_ _05504_ _05505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12182_ _00061_ clknet_leaf_77_clock u2.mem\[3\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06768__B1 _02144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06768__C2 u2.mem\[186\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11133_ _05295_ _05443_ _05461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_77_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11064_ _05390_ u2.mem\[141\]\[4\] _05412_ _05418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10015_ _04761_ _04767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_37_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07193__B1 _02556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11116__I0 _05432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12735__CLK clknet_leaf_237_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11966_ _05971_ _05980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_75_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07496__A1 _02953_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10917_ _05324_ _01054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_178_clock_I clknet_5_30_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11897_ _05940_ _01418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07113__B _02404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11419__I1 u2.mem\[163\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10848_ _05281_ _01028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12885__CLK clknet_leaf_63_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08296__I0 _03672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13567_ _01446_ clknet_leaf_15_clock u2.mem\[194\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10779_ _05240_ _01000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08996__A1 _03901_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12518_ _00397_ clknet_leaf_94_clock u2.mem\[24\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13498_ _01377_ clknet_leaf_313_clock u2.mem\[186\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_230_clock_I clknet_5_24_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12115__CLK clknet_leaf_332_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12449_ _00328_ clknet_leaf_159_clock u2.mem\[20\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09796__I0 _04609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06243__I _01553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07015__A4 _02493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07990_ u2.mem\[8\]\[15\] _03324_ _03325_ u2.mem\[4\]\[15\] _03454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12265__CLK clknet_leaf_54_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06941_ _02419_ _02420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_136_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11355__I0 _05591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08220__I0 _03568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09660_ _04543_ _04544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_5_25_0_clock_I clknet_4_12_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06872_ _02349_ _02350_ _02351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07184__B1 _02661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07723__A2 _03146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08611_ _03630_ _03542_ _03878_ _03879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_83_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09591_ _04504_ _00548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08542_ _03839_ _00164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08279__A3 _03633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08473_ _03777_ _03793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07487__B2 u2.mem\[24\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07424_ _02872_ _02877_ _02886_ _02897_ _02898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__06418__I _01918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08834__S _04015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07239__A1 u2.mem\[61\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07355_ u2.mem\[57\]\[4\] _02828_ _02829_ u2.mem\[41\]\[4\] _02830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11260__S _05536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06306_ u2.mem\[178\]\[3\] _01772_ _01773_ u2.mem\[164\]\[3\] _01810_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_332_clock clknet_5_7_0_clock clknet_leaf_332_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_136_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07286_ u2.mem\[57\]\[3\] _02554_ _02556_ u2.mem\[41\]\[3\] _02762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09025_ _04143_ _04144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06237_ _01740_ _01741_ _01742_ _01743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_1566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09787__I0 _04596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09665__S _04544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12608__CLK clknet_leaf_172_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06168_ _01638_ _01641_ _01675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07006__A4 _02484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10546__A1 _04249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_347_clock clknet_5_4_0_clock clknet_leaf_347_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07411__A1 u2.mem\[58\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06214__A2 _01582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10604__S _05131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06099_ _01578_ _01590_ _01598_ _01605_ _01606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__09464__I _04418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13190__CLK clknet_leaf_279_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07962__A2 _02503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09927_ _04614_ _04716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08211__I0 _03559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12758__CLK clknet_leaf_74_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09858_ _04670_ _00649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07714__A2 _03055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08809_ _03928_ u2.mem\[16\]\[10\] _04000_ _04003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09789_ _04599_ u2.mem\[38\]\[10\] _04628_ _04631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11820_ _05892_ _01389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11751_ _05850_ _01362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10702_ _05121_ u2.mem\[60\]\[12\] _05189_ _05190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08744__S _03963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11682_ _05798_ u2.mem\[179\]\[5\] _05800_ _05807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13421_ _01300_ clknet_leaf_297_clock u2.mem\[173\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12138__CLK clknet_leaf_38_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10633_ _05128_ u2.mem\[58\]\[15\] _05146_ _05150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13352_ _01231_ clknet_leaf_361_clock u2.mem\[162\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10564_ _05106_ u2.mem\[57\]\[5\] _05104_ _05107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11821__I1 u2.mem\[188\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12303_ _00182_ clknet_leaf_166_clock u2.mem\[11\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13283_ _01162_ clknet_leaf_360_clock u2.mem\[150\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10495_ _05064_ _00892_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12288__CLK clknet_leaf_165_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09778__I0 _04583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12234_ _00113_ clknet_leaf_52_clock u2.mem\[6\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13533__CLK clknet_leaf_318_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06205__A2 _01586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12165_ _00044_ clknet_leaf_91_clock u2.mem\[2\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06998__I _02476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10514__S _05073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09374__I _04139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06756__A3 _02223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11116_ _05432_ u2.mem\[144\]\[5\] _05444_ _05451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12096_ _01494_ clknet_leaf_214_clock u2.active_mem\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08202__I0 _03550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11047_ _05388_ u2.mem\[140\]\[3\] _05404_ _05408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08919__S _04074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09950__I0 _04700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput9 data_in_a[11] net9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11345__S _05584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12998_ _00877_ clknet_leaf_29_clock u2.mem\[54\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07469__A1 _02938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11949_ _05969_ _01441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06141__A1 _01606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08269__I0 _03575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11080__S _05422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09549__I _04144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07140_ _02618_ _02619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06444__A2 _01938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07071_ u2.mem\[60\]\[0\] _02546_ _02549_ u2.mem\[62\]\[0\] _02550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09769__I0 _04570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06022_ _01504_ _01529_ _01530_ _01531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11576__I0 _05711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12900__CLK clknet_leaf_75_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06701__I _02103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07973_ u2.mem\[61\]\[15\] _02559_ _02561_ u2.mem\[63\]\[15\] _03437_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09712_ _04576_ u2.mem\[37\]\[3\] _04567_ _04577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06924_ _02402_ _02403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_142_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07157__B1 _02634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10000__I0 _04714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09643_ _04485_ u2.mem\[35\]\[9\] _04532_ _04534_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09941__I0 _04691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06855_ u2.mem\[169\]\[5\] _02141_ _02143_ u2.mem\[147\]\[5\] _02334_ _02335_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_82_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09574_ _04493_ _00542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06786_ u2.mem\[185\]\[3\] _02120_ _02116_ u2.mem\[182\]\[3\] u2.mem\[144\]\[3\]
+ _02114_ _02268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_55_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08525_ _03828_ _00158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13406__CLK clknet_leaf_304_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08456_ _03676_ u2.mem\[8\]\[4\] _03783_ _03784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06132__A1 _01638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07475__A4 _02947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07407_ _02508_ _02881_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08387_ _03702_ u2.mem\[6\]\[10\] _03738_ _03741_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_271_clock clknet_5_20_0_clock clknet_leaf_271_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_137_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10067__I0 _04799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07338_ u2.mem\[44\]\[4\] _02654_ _02655_ u2.mem\[42\]\[4\] _02813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09621__A2 _04441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07632__A1 u2.mem\[32\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07269_ _02358_ _02745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09395__S _04376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09008_ data_in_trans\[2\].data_sync _04130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_286_clock clknet_5_20_0_clock clknet_leaf_286_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_3_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06840__C1 _02092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10280_ _04932_ _00809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_126_clock_I clknet_5_15_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12580__CLK clknet_leaf_98_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10334__S _04959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06199__A1 u2.mem\[190\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06199__B2 u2.mem\[194\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07935__A2 _02573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_0_clock clknet_5_0_0_clock clknet_leaf_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_120_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11319__I0 _05550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10133__I _04840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09932__I0 _04681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12921_ _00800_ clknet_leaf_159_clock u2.mem\[49\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11495__A2 _05690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_224_clock clknet_5_25_0_clock clknet_leaf_224_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12852_ _00731_ clknet_leaf_90_clock u2.mem\[45\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06371__A1 u2.mem\[147\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06371__B2 u2.mem\[169\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11803_ _05882_ _01382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12783_ _00662_ clknet_leaf_322_clock u2.mem\[41\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13086__CLK clknet_leaf_267_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11734_ _05839_ _05840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08474__S _03793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_239_clock clknet_5_19_0_clock clknet_leaf_239_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11665_ _05796_ u2.mem\[178\]\[4\] _05787_ _05797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06674__A2 _02156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10058__I0 _04792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13404_ _01283_ clknet_leaf_305_clock u2.mem\[170\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10616_ _05140_ _00937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11596_ _05753_ _01304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13335_ _01214_ clknet_leaf_17_clock u2.mem\[159\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06426__A2 _01924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08671__I0 _03917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10547_ _05094_ _05095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12923__CLK clknet_leaf_252_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06831__C1 u2.mem\[181\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13266_ _01145_ clknet_leaf_295_clock u2.mem\[147\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10478_ _04998_ u2.mem\[55\]\[3\] _05051_ _05055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12217_ _00096_ clknet_leaf_53_clock u2.mem\[5\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10244__S _04905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13197_ _01076_ clknet_leaf_277_clock u2.mem\[136\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07617__I _02616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07926__A2 _02531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12148_ _00027_ clknet_leaf_74_clock u2.mem\[1\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12079_ net13 clknet_2_1__leaf_clock_a data_in_trans\[15\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_328_clock_I clknet_5_7_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12303__CLK clknet_leaf_166_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06640_ _02027_ _02032_ _02125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06362__B2 u2.mem\[148\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06571_ u2.mem\[164\]\[0\] _02051_ _02055_ u2.mem\[178\]\[0\] _02056_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10297__I0 _04920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08310_ _03683_ _03684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09290_ _04256_ u2.mem\[27\]\[2\] _04313_ _04316_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06114__A1 u2.mem\[178\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06114__B2 u2.mem\[164\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08241_ _03636_ _00066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06665__A2 _02077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08172_ _03593_ _00040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07123_ _02388_ _02390_ _02484_ _02483_ _02602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_88_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06968__A3 _02446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07054_ _02532_ _02533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11549__I0 _05713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06005_ u2.driver_mem\[2\] _01513_ _01514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10154__S _04851_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10221__I0 _04893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07956_ _03416_ _03417_ _03418_ _03419_ _03420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_87_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08559__S _03846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06907_ _02385_ _02386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input28_I mem_address_a[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10888__I _05004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07887_ u2.mem\[61\]\[13\] _02559_ _02561_ u2.mem\[63\]\[13\] _03353_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09626_ _04524_ _00563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08358__I _03722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06838_ _02315_ _02316_ _02317_ _02318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06353__A1 u2.mem\[193\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09557_ _04481_ _00537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06769_ u2.mem\[164\]\[3\] _02051_ _02055_ u2.mem\[178\]\[3\] _02251_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08508_ _03816_ _00153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10288__I0 _04911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_52_clock_I clknet_5_12_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09488_ _04437_ _00512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08439_ _03772_ _00128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12946__CLK clknet_leaf_233_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09189__I _04248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11450_ _05633_ u2.mem\[165\]\[4\] _05654_ _05660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11788__I0 _05872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10401_ _03683_ _05007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06408__A2 _01887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11381_ _05587_ u2.mem\[161\]\[1\] _05616_ _05618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13120_ _00999_ clknet_leaf_244_clock u2.mem\[62\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10332_ _04918_ u2.mem\[51\]\[14\] _04959_ _04962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_277_clock_I clknet_5_21_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13051_ _00930_ clknet_leaf_254_clock u2.mem\[58\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10263_ _04922_ _04923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_127_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10212__I0 _04885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07908__A2 _03246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12002_ _00014_ clknet_leaf_42_clock u2.mem\[0\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09853__S _04666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06341__I _01843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10194_ _04804_ u2.mem\[48\]\[9\] _04875_ _04877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12326__CLK clknet_leaf_85_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11960__I0 _05911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08469__S _03788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_163_clock clknet_5_26_0_clock clknet_leaf_163_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12904_ _00783_ clknet_leaf_51_clock u2.mem\[48\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12476__CLK clknet_leaf_181_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06344__A1 u2.mem\[172\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07541__B1 _02991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06344__B2 u2.mem\[150\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12835_ _00714_ clknet_leaf_146_clock u2.mem\[44\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07105__C _02551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10279__I0 _04902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_178_clock clknet_5_30_0_clock clknet_leaf_178_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08097__A1 _03479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12766_ _00645_ clknet_leaf_203_clock u2.mem\[40\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11717_ _05828_ _01350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12697_ _00576_ clknet_leaf_111_clock u2.mem\[35\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11648_ _05758_ u2.mem\[177\]\[5\] _05778_ _05785_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_101_clock clknet_5_11_0_clock clknet_leaf_101_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_156_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput12 data_in_a[14] net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11779__I0 _05864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput23 inverter_select_a net23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput34 mem_write_n_a net34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08644__I0 _03831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11579_ _05742_ _01298_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13318_ _01197_ clknet_leaf_301_clock u2.mem\[156\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_116_clock clknet_5_14_0_clock clknet_leaf_116_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13249_ _01128_ clknet_leaf_285_clock u2.mem\[145\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07347__I _02545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10203__I0 _04813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07810_ u2.mem\[58\]\[12\] _03275_ _03276_ u2.mem\[36\]\[12\] _03277_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08572__A2 _03606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13251__CLK clknet_leaf_285_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08790_ _03992_ _00259_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09562__I _04157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07780__B1 _03100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12819__CLK clknet_leaf_60_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07741_ u2.mem\[1\]\[11\] _03028_ _03029_ u2.mem\[7\]\[11\] _03209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11703__I0 _05790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09372__I1 u2.mem\[29\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07672_ u2.mem\[29\]\[9\] _03066_ _03067_ u2.mem\[11\]\[9\] _03142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07082__I _02560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09411_ _04391_ u2.mem\[29\]\[15\] _04385_ _04392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06623_ _02022_ _02108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12969__CLK clknet_leaf_125_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09342_ _04335_ _04346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_55_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06554_ _02038_ _02039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08088__A1 _01976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08906__I _04050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09273_ _04289_ _04305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_166_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06485_ u2.mem\[0\]\[13\] _01973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11332__I _05504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08224_ _03608_ _03624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09938__S _04719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10690__I0 _05110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11993__CLK clknet_leaf_318_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08155_ _03582_ _03583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08635__I0 _03822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07106_ _02584_ _02585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08086_ data_in_trans\[14\].data_sync _03533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12349__CLK clknet_leaf_202_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07037_ _02407_ _02408_ _02498_ _02487_ _02516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_161_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06810__A2 _02156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08012__A1 _01612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10745__I1 u2.mem\[61\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11942__I0 _05222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_80_clock clknet_5_8_0_clock clknet_leaf_80_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_29_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12499__CLK clknet_leaf_123_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08988_ _04114_ _00335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07939_ _03400_ _03401_ _03402_ _03403_ _03404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_29_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09363__I1 u2.mem\[29\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10950_ _05346_ u2.mem\[134\]\[3\] _05337_ _05347_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10411__I _03696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06326__A1 u2.mem\[190\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06326__B2 u2.mem\[194\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_95_clock clknet_5_10_0_clock clknet_leaf_95_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_95_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09609_ _04514_ _00556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06877__A2 _02353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10881_ _05302_ _01040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12620_ _00499_ clknet_leaf_190_clock u2.mem\[31\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12551_ _00430_ clknet_leaf_115_clock u2.mem\[26\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06629__A2 _02002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11622__A2 _05769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11502_ _05695_ _01268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09848__S _04661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10681__I0 _05101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12482_ _00361_ clknet_leaf_164_clock u2.mem\[22\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13124__CLK clknet_leaf_23_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07841__A4 _03307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11433_ _05650_ _01244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08626__I0 _03813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_33_clock clknet_5_3_0_clock clknet_leaf_33_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11364_ _05607_ _05608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_152_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10315_ _04952_ _00824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06262__B1 _01737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13103_ _00982_ clknet_leaf_312_clock u2.mem\[61\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11295_ _05564_ _01192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07167__I _02502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13034_ _00913_ clknet_leaf_326_clock u2.mem\[56\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10246_ _04601_ _04911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08003__A1 u2.active_mem\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08003__B2 u2.active_mem\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_48_clock clknet_5_7_0_clock clknet_leaf_48_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11933__I0 _05213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11618__S _05760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10177_ _04867_ _00771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06565__A1 _02031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07762__B1 _03140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07116__B _02468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06317__A1 u2.mem\[158\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07514__B1 _02888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06317__B2 u2.mem\[151\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11353__S _05598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12818_ _00697_ clknet_leaf_147_clock u2.mem\[43\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07630__I _02447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07817__B2 u2.mem\[20\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12749_ _00628_ clknet_leaf_212_clock u2.mem\[39\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06270_ _01622_ _01775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07293__A2 _02680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08617__I0 _03804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10991__I _05372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11377__A1 _05285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07045__A2 _02521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09290__I0 _04256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06253__B1 _01658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06253__C2 u2.mem\[181\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09960_ _04735_ _00686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07077__I _02555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08911_ _04046_ u2.mem\[18\]\[14\] _04066_ _04069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12641__CLK clknet_leaf_173_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09891_ _04578_ _04691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11924__I0 _05913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08842_ _04025_ _00278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06556__A1 _02036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07753__B1 _03127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07805__I _02485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08773_ _03935_ u2.mem\[15\]\[13\] _03978_ _03980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11327__I _05499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07724_ u2.mem\[17\]\[10\] _03077_ _03078_ u2.mem\[24\]\[10\] _03193_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12791__CLK clknet_leaf_44_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08837__S _04015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06308__A1 u2.mem\[171\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06308__B2 u2.mem\[157\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_225_clock_I clknet_5_25_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07655_ u2.mem\[14\]\[9\] _03123_ _03124_ u2.mem\[12\]\[9\] _03125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06859__A2 row_select_trans\[4\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06606_ _02080_ _02015_ _02091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12021__CLK clknet_2_1__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07586_ u2.mem\[60\]\[8\] _03055_ _03056_ u2.mem\[62\]\[8\] _03057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09325_ _04246_ u2.mem\[28\]\[0\] _04336_ _04337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06537_ _02005_ _01997_ _02022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09256_ _04260_ u2.mem\[26\]\[4\] _04295_ _04296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06468_ _01927_ _01960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07284__A2 _02546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08207_ _03554_ u2.mem\[3\]\[4\] _03614_ _03615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12171__CLK clknet_leaf_209_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13297__CLK clknet_leaf_363_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09187_ _03749_ _03775_ _04247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06399_ u2.mem\[154\]\[5\] _01699_ _01701_ u2.mem\[162\]\[5\] _01900_ _01901_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__05995__I _01503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10415__I0 _05016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08138_ _03570_ u2.mem\[1\]\[11\] _03564_ _03571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08233__A1 mem_address_trans\[1\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08069_ data_in_trans\[9\].data_sync _03521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06795__A1 u2.mem\[149\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10100_ _04822_ _00739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06795__B2 u2.mem\[175\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11080_ _05428_ u2.mem\[142\]\[3\] _05422_ _05429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_1313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11915__I0 _05903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10031_ _04707_ u2.mem\[44\]\[11\] _04772_ _04776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11438__S _05646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11237__I _05528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09336__I1 u2.mem\[28\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11982_ _05225_ u2.mem\[194\]\[13\] _05985_ _05989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10933_ _05333_ _01061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11173__S _05484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10864_ _05202_ u2.mem\[129\]\[3\] _05287_ _05291_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12603_ _00482_ clknet_leaf_196_clock u2.mem\[30\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08847__I0 _04028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10795_ _05249_ _01007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12514__CLK clknet_leaf_162_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11901__S _05942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_12534_ _00413_ clknet_leaf_97_clock u2.mem\[25\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06066__I col_select_trans\[0\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07275__A2 _02495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06483__B1 _01943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12465_ _00344_ clknet_leaf_167_clock u2.mem\[21\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11700__I _05817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11416_ _05640_ _01237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07027__A2 _02503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12396_ _00275_ clknet_leaf_180_clock u2.mem\[17\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12664__CLK clknet_leaf_135_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11347_ _04417_ _05566_ _05597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06786__A1 u2.mem\[185\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07983__B1 _02598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06786__B2 u2.mem\[182\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_174_clock_I clknet_5_27_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11278_ _05513_ _05554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10229_ _04899_ _00791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13017_ _00896_ clknet_leaf_319_clock u2.mem\[55\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07735__B1 _03100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold1 output_active_trans.data_sync net45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyd_4
XFILLER_39_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09327__I1 u2.mem\[28\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07750__A3 _03216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12044__CLK clknet_leaf_299_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11083__S _05421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07440_ _02597_ _02914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10893__I0 _05294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07371_ u2.mem\[17\]\[4\] _02844_ _02845_ u2.mem\[24\]\[4\] _02846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12194__CLK clknet_leaf_238_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_99_clock_I clknet_5_10_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09110_ _03752_ _04122_ _04202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06322_ _01823_ _01824_ _01825_ _01826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07266__A2 _02457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06069__A3 _01549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09041_ _04156_ _00346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06474__B1 _01948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06253_ u2.mem\[174\]\[1\] _01656_ _01658_ u2.mem\[155\]\[1\] _01660_ u2.mem\[181\]\[1\]
+ _01759_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_148_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06184_ _01566_ _01615_ _01691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06777__A1 u2.mem\[145\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09943_ _04694_ u2.mem\[42\]\[5\] _04724_ _04726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11258__S _05537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09874_ _04679_ _00656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07726__B1 _03084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09191__A2 _04250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08825_ _04012_ _04013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_57_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08756_ _03970_ _00247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input10_I data_in_a[12] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09750__I _04566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07707_ u2.mem\[44\]\[10\] _03120_ _03121_ u2.mem\[42\]\[10\] _03176_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08687_ _03928_ u2.mem\[13\]\[10\] _03924_ _03929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12537__CLK clknet_leaf_116_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07638_ u2.mem\[16\]\[9\] _03031_ _03032_ u2.mem\[33\]\[9\] _03108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07569_ _02488_ _03040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09398__S _04376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09308_ _04274_ u2.mem\[27\]\[10\] _04323_ _04326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07257__A2 _02622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10580_ _05117_ u2.mem\[57\]\[10\] _05113_ _05118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_7_0_clock clknet_3_3_0_clock clknet_4_7_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_155_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09239_ _04284_ _00416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12250_ _00129_ clknet_leaf_57_clock u2.mem\[7\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07009__A2 _02445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06614__I _02098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11201_ _03496_ _05504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12181_ _00060_ clknet_leaf_77_clock u2.mem\[3\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06768__B2 u2.mem\[147\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11132_ _05334_ _05460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09006__I0 _04128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11063_ _05417_ _01107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12067__CLK clknet_2_1__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10014_ _04766_ _00709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13312__CLK clknet_leaf_348_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09660__I _04543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11116__I1 u2.mem\[144\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11965_ _05979_ _01447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13462__CLK clknet_leaf_346_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10916_ _05305_ u2.mem\[132\]\[4\] _05318_ _05324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08276__I _03655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07496__A2 _02958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07180__I _02527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11896_ u2.mem\[192\]\[8\] _03518_ _05937_ _05940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07113__C _02547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10847_ _05200_ u2.mem\[128\]\[2\] _05278_ _05281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10627__I0 _05121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08445__A1 _03630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13566_ _01445_ clknet_leaf_17_clock u2.mem\[194\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10778_ _05209_ u2.mem\[62\]\[6\] _05237_ _05240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06456__B1 _01947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12517_ _00396_ clknet_leaf_95_clock u2.mem\[24\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10247__S _04905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13497_ _01376_ clknet_leaf_316_clock u2.mem\[186\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12448_ _00327_ clknet_leaf_159_clock u2.mem\[20\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12379_ _00258_ clknet_leaf_207_clock u2.mem\[16\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06759__A1 u2.mem\[187\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06759__B2 u2.mem\[192\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06940_ _02389_ _02419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07708__B1 _03124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input2_I col_select_a[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09771__S _04618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11355__I1 u2.mem\[159\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06871_ col_select_trans\[5\].data_sync _01986_ _02350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11806__S _05878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08610_ _03877_ _03878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09590_ _04469_ u2.mem\[34\]\[2\] _04501_ _04504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08387__S _03738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08541_ _03804_ u2.mem\[10\]\[2\] _03836_ _03839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_5_29_0_clock_I clknet_4_14_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08472_ _03792_ _00141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10866__I0 _05204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07423_ _02889_ _02892_ _02895_ _02896_ _02897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_24_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11541__S _05708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10618__I0 _05112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07354_ _02555_ _02829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07239__A2 _02666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09011__S _04124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06305_ _01808_ _01809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_164_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07285_ u2.mem\[37\]\[3\] _02540_ _02542_ u2.mem\[59\]\[3\] _02761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09024_ data_in_trans\[5\].data_sync _04143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06236_ u2.mem\[146\]\[1\] _01692_ _01694_ u2.mem\[186\]\[1\] _01742_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08850__S _04024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06434__I _01923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11043__I0 _05384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06167_ u2.mem\[144\]\[0\] _01671_ _01673_ u2.mem\[182\]\[0\] _01674_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13335__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06098_ u2.mem\[175\]\[0\] _01602_ _01604_ u2.mem\[159\]\[0\] _01605_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09926_ _04715_ _00672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09681__S _04554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09857_ _04589_ u2.mem\[40\]\[7\] _04666_ _04670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13485__CLK clknet_leaf_289_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08808_ _04002_ _00267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10620__S _05141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09788_ _04630_ _00619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08739_ _03960_ _00240_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_122_clock_I clknet_5_15_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11750_ _05825_ u2.mem\[184\]\[0\] _05849_ _05850_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06609__I _02093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08096__I _03484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10701_ _05173_ _05189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11681_ _05806_ _01336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13420_ _01299_ clknet_leaf_298_clock u2.mem\[173\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10609__I0 _05103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10632_ _05149_ _00944_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11282__I0 _05556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13351_ _01230_ clknet_leaf_361_clock u2.mem\[162\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10563_ _05004_ _05106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06989__A1 _02410_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12302_ _00181_ clknet_leaf_181_clock u2.mem\[11\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13282_ _01161_ clknet_leaf_0_clock u2.mem\[150\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10494_ _05016_ u2.mem\[55\]\[10\] _05061_ _05064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12233_ _00112_ clknet_leaf_57_clock u2.mem\[6\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09778__I1 u2.mem\[38\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12164_ _00043_ clknet_leaf_91_clock u2.mem\[2\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_47_clock_I clknet_5_7_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11115_ _05450_ _01126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06756__A4 _02238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12095_ _01493_ clknet_leaf_214_clock u2.active_mem\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12702__CLK clknet_leaf_256_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11046_ _05407_ _01100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11626__S _05771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10530__S _05083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06913__A1 _02348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12852__CLK clknet_leaf_90_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12997_ _00876_ clknet_leaf_29_clock u2.mem\[54\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11425__I _05605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11948_ _05229_ u2.mem\[193\]\[15\] _05965_ _05969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13208__CLK clknet_leaf_281_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06141__A2 _01628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11879_ _05930_ _01410_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08269__I1 u2.mem\[4\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11273__I0 _05550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13549_ _01428_ clknet_leaf_11_clock u2.mem\[193\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_324_clock_I clknet_5_7_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12232__CLK clknet_leaf_57_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07070_ _02548_ _02549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13358__CLK clknet_leaf_356_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06021_ u2.driver_mem\[10\] _01513_ _01530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09565__I _04160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11576__I1 u2.mem\[173\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12382__CLK clknet_leaf_207_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07972_ _03420_ _03425_ _03430_ _03435_ _03436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_45_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09711_ _04575_ _04576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06923_ _02355_ _02380_ _02402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_56_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09642_ _04533_ _00570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06854_ _02331_ _02332_ _02333_ _02334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_132_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09006__S _04124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09573_ _04491_ u2.mem\[33\]\[12\] _04492_ _04493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06785_ u2.mem\[179\]\[3\] _02151_ _02153_ u2.mem\[191\]\[3\] _02267_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_1352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06380__A2 _01880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11335__I _05507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08524_ _03826_ u2.mem\[9\]\[12\] _03827_ _03828_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06429__I _01918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08455_ _03777_ _03783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_23_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06132__A2 _01576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07406_ u2.mem\[50\]\[5\] _02878_ _02879_ u2.mem\[51\]\[5\] _02880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08386_ _03740_ _00107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07880__A2 _03343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07337_ _02804_ _02805_ _02808_ _02811_ _02812_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__11070__I _05421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09676__S _04549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09209__I0 _04263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08580__S _03857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07268_ u2.mem\[16\]\[3\] _02475_ _02477_ u2.mem\[33\]\[3\] _02744_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06164__I _01670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09007_ _04129_ _00339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11016__I0 _05388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06219_ _01545_ _01555_ _01725_ _01480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06840__B1 _02078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07199_ u2.mem\[9\]\[1\] _02580_ _02582_ u2.mem\[25\]\[1\] _02677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12725__CLK clknet_leaf_72_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07396__B2 u2.mem\[30\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10414__I _03700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11319__I1 u2.mem\[157\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12875__CLK clknet_leaf_218_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09909_ _04703_ u2.mem\[41\]\[9\] _04701_ _04704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11446__S _05655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12920_ _00799_ clknet_leaf_138_clock u2.mem\[49\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07699__A2 _03031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12851_ _00730_ clknet_leaf_86_clock u2.mem\[45\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12105__CLK clknet_leaf_63_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06371__A2 _01675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_273_clock_I clknet_5_21_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11802_ _05870_ u2.mem\[187\]\[2\] _05879_ _05882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_92_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08755__S _03968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12782_ _00661_ clknet_leaf_253_clock u2.mem\[41\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11733_ _05354_ _05808_ _05839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XPHY_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06123__A2 _01629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08554__I _03835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12255__CLK clknet_leaf_217_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09448__I0 _04389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11664_ _05676_ _05796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13500__CLK clknet_leaf_317_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10058__I1 u2.mem\[45\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13403_ _01282_ clknet_leaf_309_clock u2.mem\[170\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10615_ _05110_ u2.mem\[58\]\[7\] _05136_ _05140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09073__A1 _04180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11595_ _05752_ u2.mem\[174\]\[2\] _05748_ _05753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09586__S _04501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06074__I _01580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13334_ _01213_ clknet_leaf_5_clock u2.mem\[159\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_3_4_0_clock clknet_0_clock clknet_3_4_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_10546_ _04249_ _05071_ _05094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_157_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11007__I0 _05380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06831__B1 _02034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10525__S _05078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06831__C2 _02038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13265_ _01144_ clknet_leaf_295_clock u2.mem\[147\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10477_ _05054_ _00884_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12216_ _00095_ clknet_leaf_51_clock u2.mem\[5\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13196_ _01075_ clknet_leaf_277_clock u2.mem\[136\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12147_ _00026_ clknet_leaf_73_clock u2.mem\[1\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07139__A1 _02473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12078_ data_in_trans\[14\].A clknet_leaf_343_clock data_in_trans\[14\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08187__I0 _03575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11029_ _05397_ _01093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_331_clock clknet_5_7_0_clock clknet_leaf_331_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_64_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13030__CLK clknet_leaf_32_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06570_ _02054_ _02055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_346_clock clknet_5_4_0_clock clknet_leaf_346_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_127_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08240_ _03539_ u2.mem\[4\]\[0\] _03635_ _03636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09439__I0 _04380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08464__I _03777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13180__CLK clknet_leaf_275_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08171_ _03559_ u2.mem\[2\]\[6\] _03590_ _03593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11246__I0 _05514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12748__CLK clknet_leaf_211_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07122_ _02600_ _02601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07614__A2 _03083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07053_ _02454_ _02496_ _02497_ _02411_ _02532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__06968__A4 _02393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10435__S _05030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07808__I _02494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11549__I1 u2.mem\[171\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06004_ _01512_ _01513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12898__CLK clknet_leaf_230_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06712__I _02136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07378__A1 _02843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_6_0_clock clknet_4_3_0_clock clknet_5_6_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07955_ u2.mem\[27\]\[15\] _03254_ _03255_ u2.mem\[35\]\[15\] _03419_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08178__I0 _03566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12128__CLK clknet_leaf_37_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06906_ _02364_ _02371_ _02375_ _02384_ _02385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_101_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08878__A1 _03583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08639__I _03879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07886_ _03336_ _03341_ _03346_ _03351_ _03352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_28_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09625_ _04467_ u2.mem\[35\]\[1\] _04522_ _04524_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06837_ u2.mem\[159\]\[5\] _02107_ _02109_ u2.mem\[149\]\[5\] _02317_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12278__CLK clknet_leaf_101_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09556_ _04480_ u2.mem\[33\]\[7\] _04474_ _04481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06768_ u2.mem\[169\]\[3\] _02142_ _02144_ u2.mem\[147\]\[3\] _02158_ u2.mem\[186\]\[3\]
+ _02250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_43_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13523__CLK clknet_leaf_15_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08507_ _03815_ u2.mem\[9\]\[7\] _03809_ _03816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09487_ _04389_ u2.mem\[31\]\[14\] _04434_ _04437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07302__A1 _02774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06699_ _02180_ _02181_ _02182_ _02183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08438_ _03719_ u2.mem\[7\]\[14\] _03769_ _03772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07853__A2 _03153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08369_ _03668_ u2.mem\[6\]\[2\] _03728_ _03731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11788__I1 u2.mem\[186\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10400_ _05006_ _00855_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11380_ _05617_ _01224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07605__A2 _02913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06408__A3 _01896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10331_ _04961_ _00831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10345__S _04966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10262_ _03583_ _04863_ _04922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13050_ _00929_ clknet_leaf_44_clock u2.mem\[57\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12001_ _00013_ clknet_leaf_42_clock u2.mem\[0\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10193_ _04876_ _00778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06041__A1 col_select_trans\[2\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11960__I1 u2.mem\[194\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08169__I0 _03557_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13053__CLK clknet_leaf_259_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10080__S _04802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06497__C _01911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12903_ _00782_ clknet_leaf_140_clock u2.mem\[48\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07541__A1 _01951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06344__A2 _01654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12011__D net27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12834_ _00713_ clknet_leaf_145_clock u2.mem\[44\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08485__S _03800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12765_ _00644_ clknet_leaf_204_clock u2.mem\[40\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07402__B _02745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11716_ _05825_ u2.mem\[182\]\[0\] _05827_ _05828_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08284__I _03662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12696_ _00575_ clknet_leaf_129_clock u2.mem\[35\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11647_ _05784_ _01324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput13 data_in_a[15] net13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11779__I1 u2.mem\[186\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput24 mem_address_a[0] net24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput35 output_active_a net35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08644__I1 u2.mem\[12\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11578_ _05713_ u2.mem\[173\]\[2\] _05739_ _05742_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13317_ _01196_ clknet_leaf_301_clock u2.mem\[156\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10529_ _05084_ _00906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06280__A1 u2.mem\[187\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13248_ _01127_ clknet_leaf_272_clock u2.mem\[144\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06280__B2 u2.mem\[192\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11400__I0 _05629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13179_ _01058_ clknet_leaf_275_clock u2.mem\[133\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11086__S _05421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_270_clock clknet_5_20_0_clock clknet_leaf_270_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07740_ u2.mem\[15\]\[11\] _03025_ _03026_ u2.mem\[13\]\[11\] _03208_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12420__CLK clknet_leaf_108_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11703__I1 u2.mem\[181\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13546__CLK clknet_leaf_38_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07671_ u2.mem\[26\]\[9\] _03139_ _03140_ u2.mem\[10\]\[9\] _03141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06335__A2 _01837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08580__I0 _03806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09410_ _04176_ _04391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06622_ _02044_ _02104_ _02107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_285_clock clknet_5_20_0_clock clknet_leaf_285_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09341_ _04345_ _00457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06553_ _02015_ _02037_ _02038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_169_clock_I clknet_5_27_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12570__CLK clknet_leaf_111_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06099__A1 _01578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07296__B1 _02608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09272_ _04304_ _00429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06484_ _01969_ _01970_ _01971_ _01972_ _01461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_1538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08223_ _03623_ _00061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11219__I0 _05517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08154_ _03485_ _03581_ _03582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08635__I1 u2.mem\[12\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07105_ _02577_ _02578_ _02519_ _02551_ _02584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_88_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_221_clock_I clknet_5_28_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10165__S _04856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08085_ _01973_ _03527_ _03532_ _00014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_223_clock clknet_5_25_0_clock clknet_leaf_223_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_49_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07036_ _02514_ _02515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09954__S _04729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13076__CLK clknet_leaf_24_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_29_0_clock clknet_4_14_0_clock clknet_5_29_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09753__I data_in_trans\[13\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input40_I row_select_a[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06023__A1 u2.driver_mem\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08987_ _04044_ u2.mem\[20\]\[13\] _04112_ _04114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_238_clock clknet_5_19_0_clock clknet_leaf_238_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_9_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06574__A2 _02058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07938_ u2.mem\[28\]\[14\] _03305_ _03306_ u2.mem\[31\]\[14\] _03403_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09899__I0 _04696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07869_ u2.mem\[27\]\[13\] _03254_ _03255_ u2.mem\[35\]\[13\] _03335_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06326__A2 _01702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09608_ _04487_ u2.mem\[34\]\[10\] _04511_ _04514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12913__CLK clknet_leaf_158_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10880_ _05301_ u2.mem\[130\]\[2\] _05297_ _05302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11458__I0 _05663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09539_ _04131_ _04469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08323__I0 _03693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12550_ _00429_ clknet_leaf_98_clock u2.mem\[26\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10130__I0 _04817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11501_ _05671_ u2.mem\[168\]\[2\] _05692_ _05695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12481_ _00360_ clknet_leaf_164_clock u2.mem\[22\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07039__B1 _02517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11432_ _05629_ u2.mem\[164\]\[2\] _05647_ _05650_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08626__I1 u2.mem\[12\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11630__I0 _05754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11363_ _03487_ _05606_ _05607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_125_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09864__S _04671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06262__A1 _01727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13102_ _00981_ clknet_leaf_266_clock u2.mem\[61\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10314_ _04900_ u2.mem\[51\]\[6\] _04949_ _04952_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11294_ _05554_ u2.mem\[155\]\[4\] _05558_ _05564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12006__D mem_address_trans\[0\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13033_ _00912_ clknet_leaf_328_clock u2.mem\[56\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10245_ _04910_ _00796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08003__A2 _03458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06014__A1 u2.driver_mem\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12443__CLK clknet_leaf_199_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07211__B1 _02688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11933__I1 u2.mem\[193\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10176_ _04786_ u2.mem\[48\]\[1\] _04865_ _04867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13569__CLK clknet_leaf_14_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06565__A2 _02041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07183__I _02532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11697__I0 _05798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07116__C _02551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11634__S _05770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09104__S _04197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12817_ _00696_ clknet_leaf_146_clock u2.mem\[43\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_170_clock_I clknet_5_27_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07278__B1 _02658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07132__B _02404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10121__I0 _04808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12748_ _00627_ clknet_leaf_211_clock u2.mem\[39\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08943__S _04084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12679_ _00558_ clknet_leaf_130_clock u2.mem\[34\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08617__I1 u2.mem\[12\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11377__A2 _05606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13099__CLK clknet_leaf_245_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09290__I1 u2.mem\[27\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07358__I _02564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06253__A1 u2.mem\[174\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06253__B2 u2.mem\[155\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08910_ _04068_ _00303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_30_0_clock clknet_4_15_0_clock clknet_5_30_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_48_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10713__S _05196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09890_ _04690_ _00661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_95_clock_I clknet_5_10_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11924__I1 u2.mem\[193\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08841_ _04023_ u2.mem\[17\]\[4\] _04024_ _04025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12936__CLK clknet_leaf_324_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08772_ _03979_ _00254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07723_ u2.mem\[23\]\[10\] _03146_ _03147_ u2.mem\[22\]\[10\] _03192_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07654_ _02527_ _03124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07821__I _02545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06605_ u2.mem\[151\]\[0\] _02085_ _02087_ u2.mem\[158\]\[0\] u2.mem\[193\]\[0\]
+ _02089_ _02090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07585_ _02548_ _03056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09324_ _04335_ _04336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_146_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06536_ u2.mem\[176\]\[0\] _02004_ _02014_ u2.mem\[172\]\[0\] _02020_ u2.mem\[189\]\[0\]
+ _02021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__10112__I0 _04799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09255_ _04289_ _04295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06467_ u2.mem\[192\]\[9\] _01929_ _01959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09748__I data_in_trans\[12\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08206_ _03608_ _03614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06492__A1 _01976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09186_ _04118_ _04246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06398_ _01897_ _01898_ _01899_ _01900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_leaf_162_clock clknet_5_26_0_clock clknet_leaf_162_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11612__I0 _05752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08137_ _03525_ _03570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08233__A2 mem_address_trans\[0\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06244__A1 u2.mem\[184\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12466__CLK clknet_leaf_162_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07441__B1 _02914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08068_ _01954_ _03517_ _03520_ _00009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07019_ _02410_ _02391_ _02383_ _02498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_150_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_177_clock clknet_5_27_0_clock clknet_leaf_177_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_108_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10030_ _04775_ _00716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11915__I1 u2.mem\[193\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08099__I mem_address_trans\[0\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_3_0_clock clknet_3_1_0_clock clknet_4_3_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_5_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_100_clock clknet_5_11_0_clock clknet_leaf_100_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_57_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11981_ _05988_ _01454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10932_ _05307_ u2.mem\[133\]\[5\] _05326_ _05333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08827__I _04014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10863_ _05290_ _01034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_115_clock clknet_5_14_0_clock clknet_leaf_115_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_140_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12602_ _00481_ clknet_leaf_113_clock u2.mem\[29\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10103__I0 _04790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_10794_ _05225_ u2.mem\[62\]\[13\] _05247_ _05249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12533_ _00412_ clknet_leaf_98_clock u2.mem\[25\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11851__I0 _05911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13241__CLK clknet_leaf_272_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09658__I _04440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12464_ _00343_ clknet_leaf_173_clock u2.mem\[21\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07680__B1 _03081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12809__CLK clknet_leaf_139_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11415_ _05627_ u2.mem\[163\]\[1\] _05638_ _05640_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12395_ _00274_ clknet_leaf_179_clock u2.mem\[17\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06235__A1 u2.mem\[191\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06235__B2 u2.mem\[179\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11346_ _05596_ _01211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_117_clock_I clknet_5_14_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06786__A2 _02120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12959__CLK clknet_leaf_155_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11277_ _05553_ _01185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13016_ _00895_ clknet_leaf_319_clock u2.mem\[55\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10228_ _04898_ u2.mem\[49\]\[5\] _04896_ _04899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10159_ _04855_ _00765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10590__I0 _05124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07641__I _02502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07502__A4 _02973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12339__CLK clknet_leaf_77_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09769__S _04618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07370_ _02592_ _02845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06321_ u2.mem\[159\]\[3\] _01604_ _01595_ u2.mem\[149\]\[3\] _01825_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11842__I0 _05903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09568__I _04163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09040_ _04154_ u2.mem\[21\]\[8\] _04155_ _04156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06252_ _01752_ _01755_ _01756_ _01757_ _01758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06474__A1 u2.mem\[193\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07671__B1 _03140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12489__CLK clknet_leaf_121_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06183_ u2.mem\[170\]\[0\] _01687_ _01689_ u2.mem\[156\]\[0\] _01690_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10507__I _04862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07088__I _02419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_94_clock clknet_5_10_0_clock clknet_leaf_94_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_143_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06777__A2 _02081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07974__B2 u2.mem\[62\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09942_ _04725_ _00678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07816__I _02516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09873_ _04612_ u2.mem\[40\]\[14\] _04676_ _04679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11338__I _05510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08824_ _03483_ _03540_ _03544_ _04012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_58_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07037__B _02498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08755_ _03917_ u2.mem\[15\]\[5\] _03968_ _03970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_319_clock_I clknet_5_18_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07706_ _03171_ _03172_ _03173_ _03174_ _03175_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_26_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08686_ _03701_ _03928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_32_clock clknet_5_3_0_clock clknet_leaf_32_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07551__I _02435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07637_ u2.mem\[1\]\[9\] _03028_ _03029_ u2.mem\[7\]\[9\] _03107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11073__I _05339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13264__CLK clknet_leaf_270_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09679__S _04554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07568_ _02485_ _03039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09307_ _04325_ _00443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06519_ _02003_ _02004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11833__I0 _05872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_47_clock clknet_5_7_0_clock clknet_leaf_47_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_142_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10618__S _05141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07499_ u2.mem\[32\]\[7\] _02782_ _02783_ u2.mem\[2\]\[7\] _02971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06465__A1 _01954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09238_ _04283_ u2.mem\[25\]\[14\] _04279_ _04284_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08382__I _03727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09169_ _04154_ u2.mem\[24\]\[8\] _04236_ _04237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07009__A3 _02446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11200_ _05503_ _01158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12180_ _00059_ clknet_leaf_75_clock u2.mem\[3\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06768__A2 _02142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_3_0_clock_I clknet_4_1_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11131_ _05459_ _01133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07965__B2 u2.mem\[36\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06630__I _02114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11062_ _05388_ u2.mem\[141\]\[3\] _05413_ _05417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07717__A1 _03182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10013_ _04689_ u2.mem\[44\]\[3\] _04762_ _04766_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07193__A2 _02554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08517__I0 _03822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11964_ _05915_ u2.mem\[194\]\[5\] _05975_ _05979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10915_ _05323_ _01053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07496__A3 _02963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11895_ _05939_ _01417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_43_clock_I clknet_5_6_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06077__I col_select_trans\[2\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10846_ _05280_ _01027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12631__CLK clknet_leaf_114_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13565_ _01444_ clknet_leaf_17_clock u2.mem\[194\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10528__S _05083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10777_ _05239_ _00999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09388__I _04357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06456__A1 _01945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12516_ _00395_ clknet_leaf_99_clock u2.mem\[24\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13496_ _01375_ clknet_leaf_312_clock u2.mem\[186\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12447_ _00326_ clknet_leaf_159_clock u2.mem\[20\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10327__I _04943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12781__CLK clknet_leaf_253_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12378_ _00257_ clknet_leaf_60_clock u2.mem\[15\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_268_clock_I clknet_5_22_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07956__A1 _03416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11359__S _05597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11329_ _05584_ _05585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12011__CLK clknet_2_1__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06540__I _02024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07708__A1 u2.mem\[14\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07708__B2 u2.mem\[12\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06870_ _02348_ _02349_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08668__S _03915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07184__A2 _02660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_320_clock_I clknet_5_18_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12161__CLK clknet_leaf_154_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11094__S _05435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13287__CLK clknet_leaf_364_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08540_ _03838_ _00163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08471_ _03706_ u2.mem\[8\]\[11\] _03788_ _03792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07422_ u2.mem\[43\]\[5\] _02816_ _02817_ u2.mem\[20\]\[5\] _02896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06695__A1 _02172_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07892__B1 _02575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11815__I0 _05868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07353_ _02553_ _02828_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11621__I _05768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06304_ u2.mem\[0\]\[3\] _01808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11440__A1 _04120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06715__I _02134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07284_ u2.mem\[60\]\[3\] _02546_ _02549_ u2.mem\[62\]\[3\] _02760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09023_ _04142_ _00342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10237__I _04886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06235_ u2.mem\[191\]\[1\] _01682_ _01684_ u2.mem\[179\]\[1\] _01741_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06166_ _01672_ _01673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07947__B2 u2.mem\[4\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06097_ _01603_ _01604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09925_ _04714_ u2.mem\[41\]\[14\] _04710_ _04715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11068__I _05334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12504__CLK clknet_leaf_121_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09856_ _04669_ _00648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10901__S _05309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08578__S _03857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10554__I0 _05099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09761__I data_in_trans\[15\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08807_ _03926_ u2.mem\[16\]\[9\] _04000_ _04002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09787_ _04596_ u2.mem\[38\]\[9\] _04628_ _04630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_06999_ u2.mem\[16\]\[0\] _02475_ _02477_ u2.mem\[33\]\[0\] _02478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_73_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08738_ _03937_ u2.mem\[14\]\[14\] _03957_ _03960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12654__CLK clknet_leaf_205_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08669_ _03916_ _00214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10700_ _05188_ _00973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07883__B1 _02533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11680_ _05796_ u2.mem\[179\]\[4\] _05800_ _05806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09202__S _04252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11806__I0 _05874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10609__I1 u2.mem\[58\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10631_ _05126_ u2.mem\[58\]\[14\] _05146_ _05149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06438__A1 u2.mem\[192\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13350_ _01229_ clknet_leaf_8_clock u2.mem\[161\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10562_ _05105_ _00918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12301_ _00180_ clknet_leaf_183_clock u2.mem\[11\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06989__A2 _02391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13281_ _01160_ clknet_leaf_0_clock u2.mem\[150\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10493_ _05063_ _00891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12034__CLK clknet_leaf_289_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12232_ _00111_ clknet_leaf_57_clock u2.mem\[6\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08840__I _04014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11179__S _05483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12163_ _00042_ clknet_leaf_91_clock u2.mem\[2\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06610__A1 u2.mem\[177\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06071__C1 _01577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11114_ _05430_ u2.mem\[144\]\[4\] _05444_ _05450_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06610__B2 u2.mem\[168\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12094_ _01486_ clknet_leaf_218_clock u2.active_mem\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08738__I0 _03937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12184__CLK clknet_leaf_59_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11907__S _05942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12014__D mem_address_trans\[4\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11045_ _05386_ u2.mem\[140\]\[2\] _05404_ _05407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08488__S _03800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07166__A2 _02641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06913__A2 _02350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_3_0_0_clock clknet_0_clock clknet_3_0_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_91_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12996_ _00875_ clknet_leaf_33_clock u2.mem\[54\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11947_ _05968_ _01440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07469__A3 _02940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11642__S _05779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11670__A1 _04071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11878_ u2.mem\[192\]\[0\] _03492_ _05929_ _05930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_92_1551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09112__S _04203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06141__A3 _01637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10829_ u2.mem\[63\]\[12\] _03528_ _05268_ _05269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11441__I _05654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11273__I1 u2.mem\[154\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06535__I _02019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13548_ _01427_ clknet_leaf_12_clock u2.mem\[193\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10057__I _04783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13479_ _01358_ clknet_leaf_290_clock u2.mem\[183\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06020_ u2.driver_mem\[11\] _01508_ _01529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07929__A1 _03378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06601__A1 _02023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06270__I _01622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07971_ _03431_ _03432_ _03433_ _03434_ _03435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_99_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08729__I0 _03928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09710_ _04134_ _04575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11817__S _05888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06922_ _02377_ _02401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_171_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09581__I _04176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07157__A2 _02633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12677__CLK clknet_leaf_90_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09641_ _04482_ u2.mem\[35\]\[8\] _04532_ _04533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06853_ u2.mem\[146\]\[5\] _02155_ _02157_ u2.mem\[186\]\[5\] _02333_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06365__B1 _01672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09572_ _04464_ _04492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08197__I _03608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06784_ u2.mem\[170\]\[3\] _02146_ _02148_ u2.mem\[156\]\[3\] _02266_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08523_ _03799_ _03827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_93_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06117__B1 _01623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08454_ _03782_ _00133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07405_ _02504_ _02879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08385_ _03698_ u2.mem\[6\]\[9\] _03738_ _03740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_2_0_clock clknet_4_1_0_clock clknet_5_2_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_149_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12057__CLK clknet_2_1__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07336_ u2.mem\[58\]\[4\] _02809_ _02810_ u2.mem\[36\]\[4\] _02811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07093__A1 _02451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07267_ u2.mem\[1\]\[3\] _02465_ _02471_ u2.mem\[7\]\[3\] _02743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09209__I1 u2.mem\[25\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09006_ _04128_ u2.mem\[21\]\[1\] _04124_ _04129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08660__I _03667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06840__A1 u2.mem\[165\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06218_ _01648_ _01669_ _01724_ _01725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_69_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06840__B2 u2.mem\[163\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07198_ u2.mem\[29\]\[1\] _02565_ _02570_ u2.mem\[11\]\[1\] _02676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_151_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06149_ _01561_ _01564_ _01588_ _01656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__13452__CLK clknet_leaf_342_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06180__I _01686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09908_ _04595_ _04703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09839_ _04440_ _04659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_46_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06356__B1 _01594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12850_ _00729_ clknet_leaf_150_clock u2.mem\[45\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09145__I0 _04177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_216_clock_I clknet_5_28_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11801_ _05881_ _01381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12781_ _00660_ clknet_leaf_253_clock u2.mem\[41\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_11732_ _05838_ _01355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_5_11_0_clock_I clknet_4_5_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11663_ _05795_ _01329_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09448__I1 u2.mem\[30\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13402_ _01281_ clknet_leaf_298_clock u2.mem\[170\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07608__B1 _03078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10614_ _05139_ _00936_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08771__S _03978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11594_ _05670_ _05752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13333_ _01212_ clknet_leaf_4_clock u2.mem\[159\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12009__D net26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10545_ _04986_ _05093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10806__S _05253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06831__A1 u2.mem\[155\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13264_ _01143_ clknet_leaf_270_clock u2.mem\[147\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10476_ _04995_ u2.mem\[55\]\[2\] _05051_ _05054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12215_ _00094_ clknet_leaf_53_clock u2.mem\[5\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13195_ _01074_ clknet_leaf_273_clock u2.mem\[136\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12146_ _00025_ clknet_leaf_225_clock u2.mem\[1\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12077_ net12 clknet_2_2__leaf_clock_a data_in_trans\[14\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11028_ _05384_ u2.mem\[139\]\[1\] _05395_ _05397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11191__I0 _05470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06898__A1 _02352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08946__S _04089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09136__I0 _04164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12979_ _00858_ clknet_leaf_42_clock u2.mem\[53\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13325__CLK clknet_leaf_342_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09439__I1 u2.mem\[30\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08170_ _03592_ _00039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06265__I _01614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08681__S _03924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07121_ _02547_ _02371_ _02375_ _02498_ _02600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_146_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10716__S _05196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13475__CLK clknet_leaf_295_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07052_ _02530_ _02531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06003_ u2.select_mem_row\[0\] _01510_ _01511_ _01512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07096__I _02574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_165_clock_I clknet_5_26_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11547__S _05722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07954_ u2.mem\[40\]\[15\] _03251_ _03252_ u2.mem\[30\]\[15\] _03418_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07824__I _02539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06905_ _02378_ _02382_ _02383_ _02384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_07885_ _03347_ _03348_ _03349_ _03350_ _03351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_28_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09624_ _04523_ _00562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10250__I _04886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06836_ u2.mem\[188\]\[5\] _02103_ _02105_ u2.mem\[175\]\[5\] _02316_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09127__I0 _04151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09555_ _04150_ _04480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06767_ u2.mem\[148\]\[3\] _02129_ _02131_ u2.mem\[152\]\[3\] _02248_ _02249_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_55_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11282__S _05545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08506_ _03688_ _03815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09486_ _04436_ _00511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06698_ u2.mem\[184\]\[1\] _02071_ _01993_ _02182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07302__A2 _02775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_25_0_clock clknet_4_12_0_clock clknet_5_25_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_24_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08437_ _03771_ _00127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06175__I _01681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08368_ _03730_ _00099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07319_ u2.mem\[15\]\[4\] _02792_ _02793_ u2.mem\[13\]\[4\] _02794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07066__A1 _02544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06408__A4 _01909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08299_ _03674_ _03675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10996__I0 _05343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10330_ _04916_ u2.mem\[51\]\[13\] _04959_ _04961_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12842__CLK clknet_leaf_139_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07081__A4 _02453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10261_ _04921_ _00801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10748__I0 _05220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12000_ _00012_ clknet_leaf_28_clock u2.mem\[0\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10192_ _04801_ u2.mem\[48\]\[8\] _04875_ _04876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06041__A2 col_select_trans\[3\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10361__S _04976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12992__CLK clknet_leaf_240_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09366__I0 _04360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11173__I0 _05466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10160__I _04840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12902_ _00781_ clknet_leaf_74_clock u2.mem\[48\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11873__A1 mem_address_trans\[6\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08766__S _03973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09118__I0 _04136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12222__CLK clknet_leaf_216_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13348__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12833_ _00712_ clknet_leaf_148_clock u2.mem\[44\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12764_ _00643_ clknet_leaf_203_clock u2.mem\[40\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11715_ _05826_ _05827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_43_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12695_ _00574_ clknet_leaf_110_clock u2.mem\[35\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12372__CLK clknet_leaf_80_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09597__S _04506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11646_ _05756_ u2.mem\[177\]\[4\] _05778_ _05784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07057__A1 _02450_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput14 data_in_a[1] net14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput25 mem_address_a[1] net25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11577_ _05741_ _01297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput36 row_col_select_a net36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13316_ _01195_ clknet_leaf_300_clock u2.mem\[156\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06804__A1 _02277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10528_ _05011_ u2.mem\[56\]\[8\] _05083_ _05084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08006__B1 _03459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13247_ _01126_ clknet_leaf_272_clock u2.mem\[144\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10459_ _05018_ u2.mem\[54\]\[11\] _05040_ _05044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10739__I0 _05213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11400__I1 u2.mem\[162\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13178_ _01057_ clknet_leaf_276_clock u2.mem\[133\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12129_ _01470_ clknet_leaf_35_clock u2.driver_mem\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08572__A4 _03776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07644__I _02508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07780__A2 _03099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11164__I0 _05472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11166__I _05442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10070__I _04783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07670_ _02574_ _03140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06621_ u2.mem\[188\]\[0\] _02103_ _02105_ u2.mem\[175\]\[0\] _02106_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12715__CLK clknet_leaf_252_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09340_ _04267_ u2.mem\[28\]\[7\] _04341_ _04345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06552_ _02017_ _02036_ _02037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09271_ _04276_ u2.mem\[26\]\[11\] _04300_ _04304_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_91_clock_I clknet_5_10_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06483_ u2.mem\[193\]\[12\] _01960_ _01943_ u2.mem\[194\]\[12\] _01964_ _01972_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_21_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08222_ _03570_ u2.mem\[3\]\[11\] _03619_ _03623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11219__I1 u2.mem\[150\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12865__CLK clknet_leaf_148_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07048__A1 _02407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08153_ _03481_ _03543_ _03581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_147_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10446__S _05035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10978__I0 _05335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07104_ u2.mem\[9\]\[0\] _02580_ _02582_ u2.mem\[25\]\[0\] _02583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06256__C1 u2.mem\[162\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08084_ _03531_ _03529_ _03532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07035_ _02469_ _02431_ _02433_ _02425_ _02514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_161_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07220__B2 u2.mem\[30\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08986_ _04113_ _00334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07554__I _02456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12245__CLK clknet_leaf_73_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input33_I mem_address_a[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07937_ u2.mem\[9\]\[14\] _03302_ _03303_ u2.mem\[25\]\[14\] _03402_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11076__I _05342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12112__D _01475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07868_ u2.mem\[40\]\[13\] _03251_ _03252_ u2.mem\[30\]\[13\] _03334_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09607_ _04513_ _00555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06819_ u2.mem\[154\]\[4\] _02225_ _02226_ u2.mem\[162\]\[4\] _02299_ _02300_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_28_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12395__CLK clknet_leaf_179_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07799_ u2.mem\[16\]\[12\] _03264_ _03265_ u2.mem\[33\]\[12\] _03266_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09538_ _04468_ _00531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09520__I0 _04382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09469_ _04371_ u2.mem\[31\]\[6\] _04424_ _04427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06119__B _01553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11500_ _05694_ _01267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12480_ _00359_ clknet_leaf_164_clock u2.mem\[22\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11431_ _05649_ _01243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07039__B2 u2.mem\[20\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10969__I0 _05346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_330_clock clknet_5_7_0_clock clknet_leaf_330_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11362_ _05605_ _05606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_13101_ _00980_ clknet_leaf_266_clock u2.mem\[61\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10313_ _04951_ _00823_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06262__A2 _01554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13020__CLK clknet_leaf_258_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11293_ _05563_ _01191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13032_ _00911_ clknet_leaf_328_clock u2.mem\[56\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10244_ _04909_ u2.mem\[49\]\[10\] _04905_ _04910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11394__I0 _05623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11187__S _05492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07211__A1 u2.mem\[5\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_345_clock clknet_5_5_0_clock clknet_leaf_345_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_79_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10175_ _04866_ _00770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07762__A2 _03139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13170__CLK clknet_leaf_268_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09880__S _04683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06970__B1 _02448_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11915__S _05950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12022__D mem_address_trans\[8\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11697__I1 u2.mem\[180\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07514__A2 _02887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_113_clock_I clknet_5_14_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12816_ _00695_ clknet_leaf_147_clock u2.mem\[43\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08295__I _03671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09511__I0 _04373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12888__CLK clknet_leaf_57_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07278__B2 u2.mem\[12\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07132__C _02568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12747_ _00626_ clknet_leaf_216_clock u2.mem\[39\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12678_ _00557_ clknet_leaf_89_clock u2.mem\[34\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11629_ _05774_ _01316_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10266__S _04923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06253__A2 _01656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07450__B2 u2.mem\[4\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12268__CLK clknet_leaf_185_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10337__A1 _04095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11385__I0 _05591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_38_clock_I clknet_5_6_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08840_ _04014_ _04024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07753__A2 _03126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08771_ _03932_ u2.mem\[15\]\[12\] _03978_ _03979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07722_ _03187_ _03188_ _03189_ _03190_ _03191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_2_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07653_ _02525_ _03123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06604_ _02088_ _02089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07584_ _02545_ _03055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09502__I0 _04364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09323_ _04011_ _04334_ _04335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_80_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06535_ _02019_ _02020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10112__I1 u2.mem\[46\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11560__S _05731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09254_ _04294_ _00421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06466_ u2.mem\[0\]\[9\] _01958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08205_ _03613_ _00053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09185_ _04245_ _00401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10176__S _04865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13043__CLK clknet_leaf_26_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06492__A2 _01970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06397_ u2.mem\[152\]\[5\] _01712_ _01714_ u2.mem\[148\]\[5\] _01899_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_315_clock_I clknet_5_18_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09965__S _04734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08136_ _03569_ _00028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06453__I _01918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_4_3_0_clock_I clknet_3_1_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08067_ _03518_ _03519_ _03520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09569__I0 _04489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07992__A2 _03453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07018_ _02432_ _02497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__13193__CLK clknet_leaf_274_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07744__A2 _03034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08969_ _04026_ u2.mem\[20\]\[5\] _04102_ _04104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11128__I0 _05430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11735__S _05840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11980_ _05222_ u2.mem\[194\]\[12\] _05985_ _05988_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10931_ _05332_ _01060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06704__C2 u2.mem\[192\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10862_ _05200_ u2.mem\[129\]\[2\] _05287_ _05290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09004__I _04126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12601_ _00480_ clknet_leaf_116_clock u2.mem\[29\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10793_ _05248_ _01006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12532_ _00411_ clknet_leaf_98_clock u2.mem\[25\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08843__I _03680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11851__I1 u2.mem\[190\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12463_ _00342_ clknet_leaf_172_clock u2.mem\[21\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06483__A2 _01960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11414_ _05639_ _01236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12410__CLK clknet_leaf_112_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12394_ _00273_ clknet_leaf_134_clock u2.mem\[16\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13536__CLK clknet_leaf_318_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12017__D net30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11345_ _05595_ u2.mem\[158\]\[5\] _05584_ _05596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08480__I0 _03723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07983__A2 _02596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_284_clock clknet_5_21_0_clock clknet_leaf_284_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_153_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11276_ _05552_ u2.mem\[154\]\[3\] _05546_ _05553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11367__I0 _05587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13015_ _00894_ clknet_leaf_323_clock u2.mem\[55\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10227_ _04582_ _04898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07735__A2 _03099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09980__I0 _04694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10158_ _04808_ u2.mem\[47\]\[11\] _04851_ _04855_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_299_clock clknet_5_17_0_clock clknet_leaf_299_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_94_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10089_ _04611_ _04815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07499__A1 u2.mem\[32\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_264_clock_I clknet_5_23_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_222_clock clknet_5_28_0_clock clknet_leaf_222_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_1_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06538__I _02022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08999__A1 _04121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06320_ u2.mem\[187\]\[3\] _01632_ _01635_ u2.mem\[192\]\[3\] _01824_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07120__B1 _02598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11842__I1 u2.mem\[190\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_237_clock clknet_5_19_0_clock clknet_leaf_237_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06251_ u2.mem\[175\]\[1\] _01602_ _01631_ u2.mem\[188\]\[1\] _01757_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06474__A2 _01960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07671__A1 u2.mem\[26\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07369__I _02590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09785__S _04628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12090__CLK clknet_leaf_303_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06182_ _01688_ _01689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08471__I0 _03706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12903__CLK clknet_leaf_140_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09941_ _04691_ u2.mem\[42\]\[4\] _04724_ _04725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09872_ _04678_ _00655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07726__A2 _03083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09971__I0 _04685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08823_ _03987_ _04011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07037__C _02487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08754_ _03969_ _00246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07832__I _02564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07705_ u2.mem\[58\]\[10\] _03042_ _03043_ u2.mem\[36\]\[10\] _03174_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_6_1497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08685_ _03927_ _00219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13409__CLK clknet_leaf_305_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07636_ u2.mem\[15\]\[9\] _03025_ _03026_ u2.mem\[13\]\[9\] _03106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07567_ u2.mem\[54\]\[8\] _02881_ _02882_ u2.mem\[55\]\[8\] _03038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09306_ _04272_ u2.mem\[27\]\[9\] _04323_ _04325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10097__I0 _04782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06518_ _02000_ _02002_ _02003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08663__I _03671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12433__CLK clknet_leaf_161_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07498_ u2.mem\[45\]\[7\] _02866_ _02867_ u2.mem\[34\]\[7\] _02970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_16_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11833__I1 u2.mem\[189\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13559__CLK clknet_leaf_33_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09237_ _04173_ _04283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06449_ _01878_ _01938_ _01941_ _01944_ _01469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06465__A2 _01955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09168_ _04225_ _04236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_33_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07009__A4 _02404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08119_ _03557_ u2.mem\[1\]\[5\] _03555_ _03558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12583__CLK clknet_leaf_115_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08462__I0 _03689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09099_ _04164_ u2.mem\[22\]\[11\] _04192_ _04196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11130_ _05432_ u2.mem\[145\]\[5\] _05452_ _05459_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06911__I _02389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11349__I0 _05583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11061_ _05416_ _01106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07178__B1 _02655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10012_ _04765_ _00708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_5_7_0_clock_I clknet_4_3_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11963_ _05978_ _01446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13089__CLK clknet_leaf_241_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11264__I _05499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11521__I0 _05680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10914_ _05303_ u2.mem\[132\]\[3\] _05319_ _05323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06153__A1 _01570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11894_ u2.mem\[192\]\[7\] _03515_ _05937_ _05939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07496__A4 _02968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10845_ _05198_ u2.mem\[128\]\[1\] _05278_ _05280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09669__I _04543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08573__I _03856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13564_ _01443_ clknet_leaf_18_clock u2.mem\[194\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10776_ _05207_ u2.mem\[62\]\[5\] _05237_ _05239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08445__A3 _03776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12515_ _00394_ clknet_leaf_105_clock u2.mem\[24\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06456__A2 _01938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13495_ _01374_ clknet_leaf_313_clock u2.mem\[186\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10608__I _05130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07189__I _02560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12446_ _00325_ clknet_leaf_199_clock u2.mem\[20\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06093__I _01587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12377_ _00256_ clknet_leaf_60_clock u2.mem\[15\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08453__I0 _03672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10260__I0 _04920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11328_ _04393_ _05566_ _05584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_140_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11259_ _05541_ _01179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07169__B1 _02646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07708__A2 _03123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12306__CLK clknet_leaf_166_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06977__B _02453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11760__I0 _05837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11375__S _05607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_161_clock clknet_5_26_0_clock clknet_leaf_161_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_94_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08470_ _03791_ _00140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08684__S _03924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06144__A1 _01582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12456__CLK clknet_leaf_126_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07421_ u2.mem\[49\]\[5\] _02893_ _02894_ u2.mem\[46\]\[5\] _02895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07892__B2 u2.mem\[10\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10719__S _05196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07352_ u2.mem\[37\]\[4\] _02825_ _02826_ u2.mem\[59\]\[4\] _02827_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11815__I1 u2.mem\[188\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06303_ _01769_ _01555_ _01807_ _01482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_148_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11440__A2 _05645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07283_ u2.mem\[61\]\[3\] _02666_ _02667_ u2.mem\[63\]\[3\] _02759_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10518__I _05072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07099__I _02419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09022_ _04140_ u2.mem\[21\]\[4\] _04141_ _04142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06234_ u2.mem\[170\]\[1\] _01687_ _01689_ u2.mem\[156\]\[1\] _01740_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06165_ _01665_ _01591_ _01582_ _01672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_116_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07827__I _02553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10251__I0 _04913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06096_ _01566_ _01599_ _01603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_172_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09149__A1 _04224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_114_clock clknet_5_14_0_clock clknet_leaf_114_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07048__B _02519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09924_ _04611_ _04714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09855_ _04586_ u2.mem\[40\]\[6\] _04666_ _04669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08806_ _04001_ _00266_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06998_ _02476_ _02477_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09786_ _04629_ _00618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06383__A1 u2.mem\[171\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07580__B1 _03050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_129_clock clknet_5_14_0_clock clknet_leaf_129_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08737_ _03959_ _00239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11503__I0 _05674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09321__A1 _03630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08594__S _03867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08668_ _03914_ u2.mem\[13\]\[4\] _03915_ _03916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06135__A1 _01641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13381__CLK clknet_leaf_305_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_7_clock_I clknet_5_0_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07619_ u2.mem\[39\]\[8\] _03088_ _03089_ u2.mem\[48\]\[8\] _03090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06686__A2 _02156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08599_ _03871_ _00189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07883__B2 u2.mem\[46\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11812__I _05887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12949__CLK clknet_leaf_67_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10630_ _05148_ _00943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11806__I1 u2.mem\[187\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06438__A2 _01931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10561_ _05103_ u2.mem\[57\]\[4\] _05104_ _05105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12300_ _00179_ clknet_leaf_181_clock u2.mem\[11\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06989__A3 _02424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10490__I0 _05011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13280_ _01159_ clknet_leaf_0_clock u2.mem\[150\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10492_ _05014_ u2.mem\[55\]\[9\] _05061_ _05063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12231_ _00110_ clknet_leaf_52_clock u2.mem\[6\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_212_clock_I clknet_5_29_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12162_ _00041_ clknet_leaf_153_clock u2.mem\[2\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08060__A1 _01945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12329__CLK clknet_leaf_125_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11113_ _05449_ _01125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06071__B1 _01572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06071__C2 u2.mem\[193\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12093_ _00017_ clknet_leaf_363_clock u3.enable vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06610__A2 _02092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08738__I1 u2.mem\[14\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11044_ _05406_ _01099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08363__A2 _03726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06374__A1 _01844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12479__CLK clknet_leaf_163_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12995_ _00874_ clknet_leaf_323_clock u2.mem\[54\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12030__D row_select_trans\[2\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06088__I _01594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11946_ _05227_ u2.mem\[193\]\[14\] _05965_ _05968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_93_clock clknet_5_10_0_clock clknet_leaf_93_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11670__A2 _05769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11877_ _05928_ _05929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06141__A4 _01647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10828_ _05252_ _05268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_125_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10338__I _04965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08674__I0 _03919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13547_ _01426_ clknet_leaf_35_clock u2.mem\[193\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10759_ _05228_ _00992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10481__I0 _05001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13104__CLK clknet_leaf_243_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13478_ _01357_ clknet_leaf_290_clock u2.mem\[183\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12429_ _00308_ clknet_leaf_196_clock u2.mem\[19\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07929__A2 _03383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_31_clock clknet_5_3_0_clock clknet_leaf_31_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_154_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07970_ u2.mem\[43\]\[15\] _03282_ _03283_ u2.mem\[20\]\[15\] _03434_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13254__CLK clknet_leaf_291_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06601__A2 _02033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08729__I1 u2.mem\[14\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06921_ _02374_ _02400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_68_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_46_clock clknet_5_7_0_clock clknet_leaf_46_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_95_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09640_ _04521_ _04532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_28_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06852_ u2.mem\[179\]\[5\] _02150_ _02152_ u2.mem\[191\]\[5\] _02332_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10801__I _05252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06365__A1 u2.mem\[144\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07562__B1 _03032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09571_ _04166_ _04491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06783_ _02261_ _02262_ _02263_ _02264_ _02265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_23_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08522_ _03709_ _03826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11833__S _05896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06117__A1 u2.mem\[167\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06117__B2 u2.mem\[183\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08453_ _03672_ u2.mem\[8\]\[3\] _03778_ _03782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07865__A1 _01969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_161_clock_I clknet_5_26_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07404_ _02502_ _02878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08384_ _03739_ _00106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07335_ _02499_ _02810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10472__I0 _04987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07093__A2 _02452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07266_ u2.mem\[15\]\[3\] _02457_ _02461_ u2.mem\[13\]\[3\] _02742_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09005_ _04127_ _04128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06217_ _01674_ _01697_ _01718_ _01723_ _01724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_136_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07197_ u2.mem\[26\]\[1\] _02673_ _02674_ u2.mem\[10\]\[1\] _02675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06840__A2 _02075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07557__I _02464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09973__S _04740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06148_ u2.mem\[189\]\[0\] _01650_ _01652_ u2.mem\[176\]\[0\] u2.mem\[172\]\[0\]
+ _01654_ _01655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__08042__A1 _03500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09090__I0 _04151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11079__I _05345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_5_21_0_clock clknet_4_10_0_clock clknet_5_21_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_06079_ _01584_ _01559_ _01585_ _01586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10912__S _05319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12621__CLK clknet_leaf_190_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_86_clock_I clknet_5_11_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09907_ _04702_ _00666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09838_ _04658_ _00641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06356__A1 u2.mem\[159\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06356__B2 u2.mem\[149\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09769_ _04570_ u2.mem\[38\]\[1\] _04618_ _04620_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12771__CLK clknet_leaf_90_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11800_ _05868_ u2.mem\[187\]\[1\] _05879_ _05881_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12780_ _00659_ clknet_leaf_253_clock u2.mem\[41\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_11731_ _05837_ u2.mem\[182\]\[5\] _05826_ _05838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10359__S _04976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06636__I _02120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12001__CLK clknet_leaf_42_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11662_ _05794_ u2.mem\[178\]\[3\] _05788_ _05795_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13127__CLK clknet_leaf_327_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13401_ _01280_ clknet_leaf_297_clock u2.mem\[170\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10613_ _05108_ u2.mem\[58\]\[6\] _05136_ _05139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11593_ _05751_ _01303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_5_15_0_clock_I clknet_4_7_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13332_ _01211_ clknet_leaf_8_clock u2.mem\[158\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10544_ _05092_ _00913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12151__CLK clknet_leaf_64_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06831__A2 _02029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_363_clock_I clknet_5_0_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13263_ _01142_ clknet_leaf_272_clock u2.mem\[147\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10475_ _05053_ _00883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10215__I0 _04889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09883__S _04683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12214_ _00093_ clknet_leaf_68_clock u2.mem\[5\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09081__I0 _04136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13194_ _01073_ clknet_leaf_272_clock u2.mem\[135\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12145_ _00024_ clknet_leaf_218_clock u2.mem\[1\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12025__D net37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10822__S _05263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12076_ data_in_trans\[13\].A clknet_leaf_343_clock data_in_trans\[13\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11027_ _05396_ _01092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08298__I _03506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06347__B2 u2.mem\[183\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11191__I1 u2.mem\[149\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06898__A2 _02376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11653__S _05788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12978_ _00857_ clknet_leaf_250_clock u2.mem\[53\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08895__I0 _04030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11929_ _05958_ _01432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08962__S _04097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06546__I _02006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07120_ u2.mem\[23\]\[0\] _02596_ _02598_ u2.mem\[22\]\[0\] _02599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_1494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08761__I _03962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07051_ _02413_ _02431_ _02433_ _02463_ _02530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_173_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06822__A2 _02300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06002_ _01505_ _01502_ _01511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08024__A1 _03483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10906__A1 _04095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_108_clock_I clknet_5_11_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10732__S _05205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06586__A1 _02015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07953_ u2.mem\[32\]\[15\] _03248_ _03249_ u2.mem\[2\]\[15\] _03417_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08202__S _03609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06904_ _02351_ _02383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_07884_ u2.mem\[43\]\[13\] _03282_ _03283_ u2.mem\[20\]\[13\] _03350_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06338__A1 _01814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07535__B1 _02921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09623_ _04463_ u2.mem\[35\]\[0\] _04522_ _04523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06835_ u2.mem\[187\]\[5\] _02100_ _02101_ u2.mem\[192\]\[5\] _02315_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08936__I _04073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09554_ _04479_ _00536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06766_ _02246_ _02247_ _02248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12024__CLK clknet_leaf_289_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08505_ _03814_ _00152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09485_ _04387_ u2.mem\[31\]\[13\] _04434_ _04436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08886__I0 _04021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06697_ u2.mem\[167\]\[1\] _02059_ _02061_ u2.mem\[183\]\[1\] _02181_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11362__I _05605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10693__I0 _05112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08436_ _03715_ u2.mem\[7\]\[13\] _03769_ _03771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12174__CLK clknet_leaf_210_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08367_ _03664_ u2.mem\[6\]\[1\] _03728_ _03730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07318_ _02460_ _02793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08298_ _03506_ _03674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07249_ u2.mem\[23\]\[2\] _02680_ _02681_ u2.mem\[22\]\[2\] _02726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10260_ _04920_ u2.mem\[49\]\[15\] _04914_ _04921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08015__A1 u3.data vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10191_ _04864_ _04875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_121_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07774__B1 _03092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08112__S _03546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11537__I _05676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09366__I1 u2.mem\[29\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11173__I1 u2.mem\[148\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12901_ _00780_ clknet_leaf_74_clock u2.mem\[48\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11873__A2 mem_address_trans\[7\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12832_ _00711_ clknet_leaf_145_clock u2.mem\[44\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08846__I _03684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12763_ _00642_ clknet_leaf_203_clock u2.mem\[40\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11272__I _05507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11714_ _04179_ _05808_ _05826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_42_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10684__I0 _05103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12694_ _00573_ clknet_leaf_92_clock u2.mem\[35\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11645_ _05783_ _01323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12667__CLK clknet_leaf_195_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07057__A2 _02482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput15 data_in_a[2] net15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11576_ _05711_ u2.mem\[173\]\[1\] _05739_ _05741_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput26 mem_address_a[2] net26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput37 row_select_a[0] net37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13315_ _01194_ clknet_leaf_300_clock u2.mem\[156\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06804__A2 _02282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10527_ _05072_ _05083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_122_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10458_ _05043_ _00876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13246_ _01125_ clknet_leaf_272_clock u2.mem\[144\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11648__S _05778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13177_ _01056_ clknet_leaf_275_clock u2.mem\[133\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10389_ _04997_ _04998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07765__B1 _03073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09118__S _04203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12128_ _01469_ clknet_leaf_37_clock u2.driver_mem\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12059_ net18 clknet_2_1__leaf_clock_a data_in_trans\[5\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12047__CLK clknet_2_2__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11313__A1 _05411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11164__I1 u2.mem\[147\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06985__B _02463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11383__S _05616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06620_ _02057_ _02104_ _02105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06740__A1 _02219_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06551_ _02009_ _01989_ _02036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12197__CLK clknet_leaf_72_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13442__CLK clknet_leaf_356_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09270_ _04303_ _00428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10675__I0 _05093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07296__A2 _02606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06099__A3 _01598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_34_clock_I clknet_5_3_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06482_ u2.mem\[192\]\[12\] _01929_ _01971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08221_ _03622_ _00060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08152_ _03580_ _00033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07048__A2 _02408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07103_ _02581_ _02582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06256__B1 _01698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06256__C2 _01700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08083_ data_in_trans\[13\].data_sync _03531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_3_0_clock_I clknet_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07034_ _02490_ _02501_ _02506_ _02512_ _02513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_66_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_259_clock_I clknet_5_23_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10462__S _05045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07835__I _02579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08985_ _04041_ u2.mem\[20\]\[12\] _04112_ _04113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07936_ u2.mem\[29\]\[14\] _03299_ _03300_ u2.mem\[11\]\[14\] _03401_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08867__S _04042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input26_I mem_address_a[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07867_ u2.mem\[32\]\[13\] _03248_ _03249_ u2.mem\[2\]\[13\] _03333_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_311_clock_I clknet_5_17_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09606_ _04485_ u2.mem\[34\]\[9\] _04511_ _04513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08666__I _03675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06818_ _02296_ _02297_ _02298_ _02299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07798_ _02476_ _03265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09537_ _04467_ u2.mem\[33\]\[1\] _04465_ _04468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06749_ u2.mem\[185\]\[2\] _02121_ _02123_ u2.mem\[173\]\[2\] _02232_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_145_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10666__I0 _05124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09520__I1 u2.mem\[32\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09468_ _04426_ _00503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08419_ _03761_ _00119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10637__S _05152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09399_ _04383_ _00477_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10418__I0 _05018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07039__A2 _02515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11430_ _05627_ u2.mem\[164\]\[1\] _05647_ _05649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10043__A1 _03904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11361_ _04439_ _05274_ _05605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_4_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06798__B2 u2.mem\[183\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13100_ _00979_ clknet_leaf_264_clock u2.mem\[61\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10312_ _04898_ u2.mem\[51\]\[5\] _04949_ _04951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11292_ _05552_ u2.mem\[155\]\[3\] _05559_ _05563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10243_ _04598_ _04909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13031_ _00910_ clknet_leaf_326_clock u2.mem\[56\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11543__A1 _04310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07747__B1 _03115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11394__I1 u2.mem\[162\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10174_ _04782_ u2.mem\[48\]\[0\] _04865_ _04866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07211__A2 _02687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13315__CLK clknet_leaf_300_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10171__I _04862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08777__S _03978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06970__B2 u2.mem\[34\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13465__CLK clknet_leaf_346_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06722__A1 u2.mem\[164\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06722__B2 u2.mem\[178\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12815_ _00694_ clknet_leaf_146_clock u2.mem\[43\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10657__I0 _05115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09511__I1 u2.mem\[32\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07278__A2 _02657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12746_ _00625_ clknet_leaf_50_clock u2.mem\[38\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12677_ _00556_ clknet_leaf_90_clock u2.mem\[34\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11730__I _03679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10409__I0 _05011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11628_ _05752_ u2.mem\[176\]\[2\] _05771_ _05774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06238__B1 _01680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11559_ _05730_ _05731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06789__A1 _02255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09027__I0 _04145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_260_clock_I clknet_5_23_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10282__S _04933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13229_ _01108_ clknet_leaf_286_clock u2.mem\[141\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10337__A2 _04964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07738__B1 _03022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11385__I1 u2.mem\[161\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08770_ _03962_ _03978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_97_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08687__S _03924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06961__A1 _02348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07721_ u2.mem\[28\]\[10\] _03072_ _03073_ u2.mem\[31\]\[10\] _03190_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_4_10_0_clock_I clknet_3_5_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07652_ u2.mem\[44\]\[9\] _03120_ _03121_ u2.mem\[42\]\[9\] _03122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06713__A1 u2.mem\[153\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12832__CLK clknet_leaf_145_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06603_ _01992_ _02080_ _02088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_168_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07583_ u2.mem\[61\]\[8\] _02899_ _02900_ u2.mem\[63\]\[8\] _03054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06534_ _02015_ _02018_ _02019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09322_ _04333_ _04334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10648__I0 _05106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09253_ _04258_ u2.mem\[26\]\[3\] _04290_ _04294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06465_ _01954_ _01955_ _01956_ _01957_ _01472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10457__S _05040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12982__CLK clknet_leaf_31_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08204_ _03552_ u2.mem\[3\]\[3\] _03609_ _03613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09184_ _04177_ u2.mem\[24\]\[15\] _04241_ _04245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06396_ u2.mem\[153\]\[5\] _01707_ _01709_ u2.mem\[160\]\[5\] _01898_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08135_ _03568_ u2.mem\[1\]\[10\] _03564_ _03569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06229__B1 _01734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12212__CLK clknet_leaf_67_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08066_ _03493_ _03519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07441__A2 _02913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13338__CLK clknet_leaf_9_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07017_ _02430_ _02496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__10192__S _04875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07992__A3 _03454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07729__B1 _03089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_7_0_clock_I clknet_3_3_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13488__CLK clknet_leaf_298_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06401__B1 _01721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08968_ _04103_ _00326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11128__I1 u2.mem\[145\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07919_ u2.mem\[50\]\[14\] _02503_ _02505_ u2.mem\[51\]\[14\] _03384_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_5_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08899_ _04062_ _00298_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10930_ _05305_ u2.mem\[133\]\[4\] _05326_ _05332_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06909__I _02387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06704__A1 u2.mem\[188\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06704__B2 u2.mem\[187\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10861_ _05289_ _01033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12600_ _00479_ clknet_leaf_117_clock u2.mem\[29\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_1540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10639__I0 _05097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10792_ _05222_ u2.mem\[62\]\[12\] _05247_ _05248_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_12531_ _00410_ clknet_leaf_103_clock u2.mem\[25\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12462_ _00341_ clknet_leaf_191_clock u2.mem\[21\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06644__I _02128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07680__A2 _03080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09020__I _04139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11413_ _05623_ u2.mem\[163\]\[0\] _05638_ _05639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12393_ _00272_ clknet_leaf_132_clock u2.mem\[16\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07968__B1 _02528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11344_ _05516_ _05595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12705__CLK clknet_leaf_238_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11275_ _05510_ _05552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13014_ _00893_ clknet_leaf_28_clock u2.mem\[55\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10226_ _04897_ _00790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12033__D net41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11926__S _05955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10157_ _04854_ _00764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12855__CLK clknet_leaf_133_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10088_ _04814_ _00735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_207_clock_I clknet_5_29_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09496__I0 _04356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06459__B1 _01948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12729_ _00608_ clknet_leaf_44_clock u2.mem\[37\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11460__I _03496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06250_ u2.mem\[187\]\[1\] _01633_ _01636_ u2.mem\[192\]\[1\] _01756_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12235__CLK clknet_leaf_211_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06554__I _02038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07671__A2 _03139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06181_ _01566_ _01629_ _01688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_156_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12385__CLK clknet_leaf_223_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09940_ _04718_ _04724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_104_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09871_ _04609_ u2.mem\[40\]\[13\] _04676_ _04678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07187__A1 _02639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08822_ _03656_ _04010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08753_ _03914_ u2.mem\[15\]\[4\] _03968_ _03969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07704_ u2.mem\[53\]\[10\] _03039_ _03040_ u2.mem\[56\]\[10\] _03173_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08684_ _03926_ u2.mem\[13\]\[9\] _03924_ _03927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07635_ _03101_ _03102_ _03103_ _03104_ _03105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_1908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13010__CLK clknet_leaf_237_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06162__A2 _01662_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09487__I0 _04389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07566_ u2.mem\[50\]\[8\] _02878_ _02879_ u2.mem\[51\]\[8\] _03037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09305_ _04324_ _00442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11294__I0 _05554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06517_ _01991_ _02001_ _02002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_344_clock clknet_5_5_0_clock clknet_leaf_344_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_110_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07497_ _01945_ _02780_ _02948_ _02969_ _01498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_70_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09236_ _04282_ _00415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08880__S _04051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06448_ u2.mem\[193\]\[5\] _01942_ _01943_ u2.mem\[194\]\[5\] _01934_ _01944_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_107_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13160__CLK clknet_leaf_276_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12118__D _01481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09167_ _04235_ _00393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06379_ u2.mem\[180\]\[5\] _01664_ _01667_ u2.mem\[150\]\[5\] _01881_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12728__CLK clknet_leaf_54_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09775__I _04617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_359_clock clknet_5_1_0_clock clknet_leaf_359_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08118_ _03511_ _03557_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08611__A1 _03630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06217__A3 _01718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09098_ _04195_ _00364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08049_ data_in_trans\[4\].data_sync _03506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_3_clock_I clknet_5_0_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11349__I1 u2.mem\[159\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_156_clock_I clknet_5_26_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11060_ _05386_ u2.mem\[141\]\[2\] _05413_ _05416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09411__I0 _04391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10011_ _04687_ u2.mem\[44\]\[2\] _04762_ _04765_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10650__S _05157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06925__A1 _02401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06386__C1 u2.mem\[163\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12108__CLK clknet_leaf_135_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11962_ _05913_ u2.mem\[194\]\[4\] _05975_ _05978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09015__I _04135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10913_ _05322_ _01052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11893_ _05938_ _01416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09478__I0 _04380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12258__CLK clknet_leaf_228_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10844_ _05279_ _01026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_16_0_clock clknet_4_8_0_clock clknet_5_16_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__13503__CLK clknet_leaf_331_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10097__S _04820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13563_ _01442_ clknet_leaf_16_clock u2.mem\[194\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10775_ _05238_ _00998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12514_ _00393_ clknet_leaf_162_clock u2.mem\[24\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09886__S _04683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13494_ _01373_ clknet_leaf_295_clock u2.mem\[185\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12445_ _00324_ clknet_leaf_198_clock u2.mem\[20\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12028__D row_select_trans\[1\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09650__I0 _04491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12376_ _00255_ clknet_leaf_131_clock u2.mem\[15\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11327_ _05499_ _05583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09402__I0 _04384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11258_ _05511_ u2.mem\[153\]\[3\] _05537_ _05541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11656__S _05788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10209_ _04564_ _04885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06377__C1 u2.mem\[172\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11189_ _05468_ u2.mem\[149\]\[3\] _05492_ _05496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06977__C _02455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11760__I1 u2.mem\[184\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13033__CLK clknet_leaf_328_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_358_clock_I clknet_5_1_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06144__A2 _01634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07420_ _02532_ _02894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07892__A2 _02573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09469__I0 _04371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11276__I0 _05552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07351_ _02541_ _02826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09796__S _04633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06302_ _01780_ _01784_ _01793_ _01806_ _01807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_07282_ _02741_ _02747_ _02752_ _02757_ _02758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_143_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09021_ _04123_ _04141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11028__I0 _05384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06233_ u2.mem\[173\]\[1\] _01720_ _01722_ u2.mem\[185\]\[1\] _01739_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06852__B1 _02152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10735__S _05205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06164_ _01670_ _01671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09641__I0 _04482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10251__I1 u2.mem\[49\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06095_ _01601_ _01602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09923_ _04713_ _00671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07048__C _02454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11566__S _05731_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09854_ _04668_ _00647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07843__I _02590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08805_ _03923_ u2.mem\[16\]\[8\] _04000_ _04001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09785_ _04592_ u2.mem\[38\]\[8\] _04628_ _04629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_06997_ _02429_ _02445_ _02446_ _02463_ _02476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_85_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06383__A2 _01610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07580__B2 u2.mem\[20\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08736_ _03935_ u2.mem\[14\]\[13\] _03957_ _03959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11503__I1 u2.mem\[168\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13526__CLK clknet_leaf_314_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08667_ _03905_ _03915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06135__A2 _01596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08380__I0 _03689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07618_ _02618_ _03089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08598_ _03824_ u2.mem\[11\]\[11\] _03867_ _03871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07883__A2 _02531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_283_clock clknet_5_21_0_clock clknet_leaf_283_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11267__I0 _05544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07549_ u2.mem\[40\]\[8\] _03018_ _03019_ u2.mem\[30\]\[8\] _03020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_82_clock_I clknet_5_9_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12550__CLK clknet_leaf_98_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08132__I0 _03566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06194__I _01700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07635__A2 _03102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10560_ _05094_ _05104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_167_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09880__I0 _04681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09219_ _04269_ u2.mem\[25\]\[8\] _04270_ _04271_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_298_clock clknet_5_17_0_clock clknet_leaf_298_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_148_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10491_ _05062_ _00890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12230_ _00109_ clknet_leaf_69_clock u2.mem\[6\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06922__I _02377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09632__I0 _04473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12161_ _00040_ clknet_leaf_154_clock u2.mem\[2\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_221_clock clknet_5_28_0_clock clknet_leaf_221_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06071__A1 u2.mem\[158\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11112_ _05428_ u2.mem\[144\]\[3\] _05445_ _05449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06071__B2 u2.mem\[151\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12092_ inverter_select_trans.A clknet_leaf_302_clock inverter_select_trans.data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13056__CLK clknet_leaf_243_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11043_ _05384_ u2.mem\[140\]\[1\] _05404_ _05406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08849__I _03688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08363__A3 _03633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_236_clock clknet_5_19_0_clock clknet_leaf_236_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11275__I _05510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12080__CLK clknet_leaf_303_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12994_ _00873_ clknet_leaf_236_clock u2.mem\[54\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11945_ _05967_ _01439_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08371__I0 _03672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06677__A3 _02140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11876_ _05927_ _05928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10827_ _05267_ _01021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13546_ _01425_ clknet_leaf_38_clock u2.mem\[192\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10758_ _05227_ u2.mem\[61\]\[14\] _05223_ _05228_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09871__I0 _04609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13477_ _01356_ clknet_leaf_298_clock u2.mem\[183\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10689_ _05182_ _00968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12428_ _00307_ clknet_leaf_180_clock u2.mem\[19\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09623__I0 _04463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07929__A3 _03388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11430__I0 _05627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12359_ _00238_ clknet_leaf_133_clock u2.mem\[14\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06598__C1 u2.mem\[145\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06920_ _02370_ _02399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_84_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07663__I _02560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12423__CLK clknet_leaf_128_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07011__B1 _02489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06851_ u2.mem\[170\]\[5\] _02145_ _02147_ u2.mem\[156\]\[5\] _02331_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06365__A2 _01670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07562__B2 u2.mem\[33\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09570_ _04490_ _00541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06782_ u2.mem\[176\]\[3\] _02003_ _02019_ u2.mem\[189\]\[3\] _02264_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08521_ _03825_ _00157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11497__I0 _05663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06117__A2 _01622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12573__CLK clknet_leaf_187_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_104_clock_I clknet_5_11_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08452_ _03781_ _00132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07865__A2 _03246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07403_ _02873_ _02874_ _02875_ _02876_ _02877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08383_ _03693_ u2.mem\[6\]\[8\] _03738_ _03739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07078__B1 _02556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07334_ _02494_ _02809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09862__I0 _04596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07265_ _02737_ _02738_ _02739_ _02740_ _02741_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07838__I _02584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09004_ _04126_ _04127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06216_ u2.mem\[173\]\[0\] _01720_ _01722_ u2.mem\[185\]\[0\] _01723_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06742__I _02126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07196_ _02574_ _02674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13079__CLK clknet_leaf_43_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11421__I0 _05633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06147_ _01653_ _01654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09090__I1 u2.mem\[22\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07250__B1 _02593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06078_ _01573_ _01574_ _01585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11296__S _05558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_29_clock_I clknet_5_3_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09906_ _04700_ u2.mem\[41\]\[8\] _04701_ _04702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09837_ _04615_ u2.mem\[39\]\[15\] _04654_ _04658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06356__A2 _01603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12916__CLK clknet_leaf_60_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09768_ _04619_ _00610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08719_ _03949_ _00231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11488__I0 _05674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09699_ _04566_ _04567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_54_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11730_ _03679_ _05837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06917__I _02395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11661_ _05673_ _05794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13400_ _01279_ clknet_leaf_301_clock u2.mem\[170\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10612_ _05138_ _00935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07608__A2 _03077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09853__I0 _04583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11592_ _05750_ u2.mem\[174\]\[1\] _05748_ _05751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13331_ _01210_ clknet_leaf_353_clock u2.mem\[158\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10543_ _05027_ u2.mem\[56\]\[15\] _05088_ _05092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_306_clock_I clknet_5_16_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13262_ _01141_ clknet_leaf_271_clock u2.mem\[147\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10474_ _04992_ u2.mem\[55\]\[1\] _05051_ _05053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_160_clock clknet_5_26_0_clock clknet_leaf_160_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_108_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12213_ _00092_ clknet_leaf_68_clock u2.mem\[5\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_5_19_0_clock_I clknet_4_9_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13193_ _01072_ clknet_leaf_274_clock u2.mem\[135\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12446__CLK clknet_leaf_199_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12144_ _00023_ clknet_leaf_226_clock u2.mem\[1\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07241__B1 _02542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12075_ net11 clknet_2_2__leaf_clock_a data_in_trans\[13\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_175_clock clknet_5_27_0_clock clknet_leaf_175_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_89_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07139__A4 _02384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11026_ _05380_ u2.mem\[139\]\[0\] _05395_ _05396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_46_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08592__I0 _03817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12977_ _00856_ clknet_leaf_250_clock u2.mem\[53\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08344__I0 _03710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11928_ _05209_ u2.mem\[193\]\[6\] _05955_ _05958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11859_ _04416_ _05886_ _05917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_53_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_113_clock clknet_5_14_0_clock clknet_leaf_113_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_18_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09844__I0 _04570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13529_ _01408_ clknet_leaf_316_clock u2.mem\[191\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13221__CLK clknet_leaf_281_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07050_ u2.mem\[14\]\[0\] _02526_ _02528_ u2.mem\[12\]\[0\] _02529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_12_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_128_clock clknet_5_14_0_clock clknet_leaf_128_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06822__A3 _02301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06001_ _01502_ _01510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_127_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11403__I0 _05631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08024__A2 _03484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07378__A4 _02852_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13371__CLK clknet_leaf_357_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07783__A1 u2.mem\[32\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_30_clock_I clknet_5_3_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06586__A2 _02070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07952_ u2.mem\[45\]\[15\] _02444_ _02448_ u2.mem\[34\]\[15\] _03416_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12939__CLK clknet_leaf_251_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07393__I _02447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06903_ _02381_ _02382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_07883_ u2.mem\[49\]\[13\] _02531_ _02533_ u2.mem\[46\]\[13\] _03349_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07535__A1 u2.mem\[5\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08583__I0 _03808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09622_ _04521_ _04522_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_112_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06834_ _02310_ _02311_ _02312_ _02313_ _02314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_95_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10390__I0 _04998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09553_ _04478_ u2.mem\[33\]\[6\] _04474_ _04479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06765_ u2.mem\[153\]\[3\] _02196_ _02200_ u2.mem\[160\]\[3\] _02247_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08504_ _03813_ u2.mem\[9\]\[6\] _03809_ _03814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07299__B1 _02619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_255_clock_I clknet_5_23_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09484_ _04435_ _00510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06696_ u2.mem\[164\]\[1\] _02050_ _02054_ u2.mem\[178\]\[1\] _02180_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08435_ _03770_ _00126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12319__CLK clknet_leaf_157_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08366_ _03729_ _00098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09835__I0 _04612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07317_ _02456_ _02792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11642__I0 _05752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08297_ _03673_ _00085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07568__I _02485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06274__A1 u2.mem\[184\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12469__CLK clknet_leaf_106_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07248_ _02721_ _02722_ _02723_ _02724_ _02725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_125_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07471__B1 _02891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07179_ _02525_ _02657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07223__B1 _02461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_92_clock clknet_5_10_0_clock clknet_leaf_92_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10190_ _04874_ _00777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07774__B2 u2.mem\[4\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08574__I0 _03798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12900_ _00779_ clknet_leaf_75_clock u2.mem\[48\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11754__S _05849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12831_ _00710_ clknet_leaf_149_clock u2.mem\[44\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12762_ _00641_ clknet_5_13_0_clock u2.mem\[39\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_30_clock clknet_5_3_0_clock clknet_leaf_30_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11713_ _03655_ _05825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12693_ _00572_ clknet_leaf_92_clock u2.mem\[35\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13244__CLK clknet_leaf_291_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09958__I _04718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08862__I _03705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11644_ _05754_ u2.mem\[177\]\[3\] _05779_ _05783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09826__I0 _04599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_45_clock clknet_5_6_0_clock clknet_leaf_45_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07057__A3 _02513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11575_ _05740_ _01296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput16 data_in_a[3] net16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput27 mem_address_a[3] net27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_5_30_0_clock_I clknet_4_15_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13314_ _01193_ clknet_leaf_349_clock u2.mem\[155\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput38 row_select_a[1] net38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10526_ _05082_ _00905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06804__A3 _02283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13245_ _01124_ clknet_leaf_285_clock u2.mem\[144\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12036__D row_select_trans\[5\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08006__A2 _03458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10457_ _05016_ u2.mem\[54\]\[10\] _05040_ _05043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07214__B1 _02624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13176_ _01055_ clknet_leaf_269_clock u2.mem\[132\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10388_ _04134_ _04997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07765__B2 u2.mem\[31\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12127_ _01468_ clknet_leaf_36_clock u2.driver_mem\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08102__I _03545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12058_ data_in_trans\[4\].A clknet_leaf_300_clock data_in_trans\[4\].data_sync vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07517__B2 u2.mem\[20\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11009_ _05339_ _05384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10372__I0 _04920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09134__S _04213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06985__C _02398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08317__I0 _03689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06550_ _02034_ _02035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10124__I0 _04810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06481_ _01920_ _01970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06099__A4 _01605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09868__I _04660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08220_ _03568_ u2.mem\[3\]\[10\] _03619_ _03622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09817__I0 _04586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12611__CLK clknet_leaf_94_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08151_ _03579_ u2.mem\[1\]\[15\] _03573_ _03580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11624__I0 _05746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07102_ _02418_ _02420_ _02552_ _02426_ _02581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__06256__A1 u2.mem\[148\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06256__B2 u2.mem\[154\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08082_ _01969_ _03527_ _03530_ _00013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_173_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07033_ u2.mem\[54\]\[0\] _02509_ _02511_ u2.mem\[55\]\[0\] _02512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12761__CLK clknet_leaf_141_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07205__B1 _02593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_7_0_clock_I clknet_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08213__S _03614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07756__A1 _03207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08984_ _04096_ _04112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_102_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13117__CLK clknet_leaf_261_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07935_ u2.mem\[26\]\[14\] _02573_ _02575_ u2.mem\[10\]\[14\] _03400_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07508__A1 _02975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11574__S _05739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07866_ u2.mem\[45\]\[13\] _02444_ _02448_ u2.mem\[34\]\[13\] _03332_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10363__I0 _04911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09044__S _04155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09605_ _04512_ _00554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input19_I data_in_a[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06817_ u2.mem\[148\]\[4\] _02129_ _02131_ u2.mem\[152\]\[4\] _02298_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07797_ _02474_ _03264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12141__CLK clknet_leaf_211_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06731__A2 _02211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13267__CLK clknet_leaf_5_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09536_ _04127_ _04467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10115__I0 _04801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06748_ u2.mem\[154\]\[2\] _02225_ _02226_ u2.mem\[162\]\[2\] _02230_ _02231_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_58_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09467_ _04369_ u2.mem\[31\]\[5\] _04424_ _04426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11863__I0 _05907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10918__S _05318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06679_ _01545_ _01996_ _02163_ _01474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08418_ _03681_ u2.mem\[7\]\[5\] _03759_ _03761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12291__CLK clknet_leaf_103_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07692__B1 _03100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09398_ _04382_ u2.mem\[29\]\[11\] _04376_ _04383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09808__I0 _04573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08349_ _03715_ u2.mem\[5\]\[13\] _03711_ _03716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10043__A2 _04760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11360_ _05604_ _01217_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10311_ _04950_ _00822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11291_ _05562_ _01190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09219__S _04270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13030_ _00909_ clknet_leaf_32_clock u2.mem\[56\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10242_ _04908_ _00795_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11543__A2 _05690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10452__I _05029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10173_ _04864_ _04865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_65_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09018__I data_in_trans\[4\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11484__S _05683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06970__A2 _02444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10354__I0 _04902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06707__C1 u2.mem\[181\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06183__B1 _01689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12814_ _00693_ clknet_leaf_220_clock u2.mem\[43\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09889__S _04683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10106__I0 _04792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08793__S _03990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12634__CLK clknet_leaf_114_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12745_ _00624_ clknet_leaf_53_clock u2.mem\[38\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11854__I0 _05913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12676_ _00555_ clknet_leaf_90_clock u2.mem\[34\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11627_ _05773_ _01315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12784__CLK clknet_leaf_321_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06238__A1 u2.mem\[147\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11558_ _04333_ _05729_ _05730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07986__A1 u2.mem\[18\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07001__I _02479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06789__A2 _02260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11659__S _05788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10509_ _05072_ _05073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_171_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_203_clock_I clknet_5_29_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09027__I1 u2.mem\[21\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11489_ _05687_ _01263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12014__CLK clknet_leaf_289_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11909__I1 _03533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13228_ _01107_ clknet_leaf_280_clock u2.mem\[141\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13159_ _01038_ clknet_leaf_274_clock u2.mem\[130\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10593__I0 _05126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12164__CLK clknet_leaf_91_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06961__A2 _02423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11394__S _05625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07720_ u2.mem\[9\]\[10\] _03069_ _03070_ u2.mem\[25\]\[10\] _03189_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10345__I0 _04893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07651_ _02522_ _03121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07910__A1 u2.mem\[32\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06602_ _02086_ _02087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07582_ _03024_ _03036_ _03045_ _03052_ _03053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_59_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09321_ _03630_ _03540_ _03878_ _04333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA_clkbuf_4_14_0_clock_I clknet_3_7_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06533_ _02017_ _02011_ _02018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11845__I0 _05907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09252_ _04293_ _00420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07674__B1 _03073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06464_ u2.mem\[193\]\[8\] _01942_ _01943_ u2.mem\[194\]\[8\] _01949_ _01957_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_72_1540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08203_ _03612_ _00052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_2_1__f_clock_a_I clknet_0_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09183_ _04244_ _00400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09415__A1 _04394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06395_ u2.mem\[190\]\[5\] _01702_ _01704_ u2.mem\[194\]\[5\] _01897_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06229__A1 u2.mem\[145\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08134_ _03523_ _03568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06229__B2 u2.mem\[177\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07977__A1 _03437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10820__I1 _03518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08065_ data_in_trans\[8\].data_sync _03518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07846__I _02600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07016_ _02494_ _02495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08777__I0 _03939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12507__CLK clknet_leaf_179_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10272__I _04922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06401__B2 u2.mem\[185\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08967_ _04023_ u2.mem\[20\]\[4\] _04102_ _04103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07918_ _03379_ _03380_ _03381_ _03382_ _03383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_40_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08898_ _04032_ u2.mem\[18\]\[8\] _04061_ _04062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12657__CLK clknet_leaf_224_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07849_ _02605_ _03316_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07901__A1 _03363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10860_ _05198_ u2.mem\[129\]\[1\] _05287_ _05289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09519_ _04456_ _00524_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_152_clock_I clknet_5_25_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10648__S _05157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10791_ _05231_ _05247_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12530_ _00409_ clknet_leaf_166_clock u2.mem\[25\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07665__B1 _03056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_12461_ _00340_ clknet_leaf_196_clock u2.mem\[21\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11412_ _05637_ _05638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12037__CLK clknet_2_0__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12392_ _00271_ clknet_leaf_133_clock u2.mem\[16\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07968__A1 u2.mem\[14\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07968__B2 u2.mem\[12\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11343_ _05594_ _01210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10811__I1 _03507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11274_ _05551_ _01184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12187__CLK clknet_leaf_251_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11278__I _05513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08768__I0 _03930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13013_ _00892_ clknet_leaf_29_clock u2.mem\[55\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10225_ _04895_ u2.mem\[49\]\[4\] _04896_ _04897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10182__I _04864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_5_12_0_clock clknet_4_6_0_clock clknet_5_12_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_95_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_77_clock_I clknet_5_8_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10156_ _04806_ u2.mem\[47\]\[10\] _04851_ _04854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10087_ _04813_ u2.mem\[45\]\[13\] _04811_ _04814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09193__I0 _04246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11942__S _05965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11827__I0 _05864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10989_ _05371_ _01079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12728_ _00607_ clknet_leaf_54_clock u2.mem\[37\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09211__I _04147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07120__A2 _02596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12659_ _00538_ clknet_leaf_81_clock u2.mem\[33\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06180_ _01686_ _01687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11389__S _05615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10293__S _04938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_354_clock_I clknet_5_1_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10802__I1 _03492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06631__A1 _02000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08759__I0 _03921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09870_ _04677_ _00654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08821_ _04009_ _00273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06395__B1 _01704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08752_ _03962_ _03968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_113_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08497__I _03799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09184__I0 _04177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07703_ u2.mem\[54\]\[10\] _03114_ _03115_ u2.mem\[55\]\[10\] _03172_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_6_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08683_ _03697_ _03926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07634_ u2.mem\[27\]\[9\] _03021_ _03022_ u2.mem\[35\]\[9\] _03104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06698__A1 u2.mem\[184\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07565_ _03027_ _03030_ _03033_ _03035_ _03036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_53_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10468__S _05045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09304_ _04269_ u2.mem\[27\]\[8\] _04323_ _04324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06516_ _01985_ _01986_ _02001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_167_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07647__B1 _03040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11294__I1 u2.mem\[155\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07496_ _02953_ _02958_ _02963_ _02968_ _02969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_107_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13305__CLK clknet_leaf_358_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09235_ _04281_ u2.mem\[25\]\[13\] _04279_ _04282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06447_ _01923_ _01943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09166_ _04151_ u2.mem\[24\]\[7\] _04231_ _04235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06378_ u2.mem\[174\]\[5\] _01657_ _01659_ u2.mem\[155\]\[5\] _01661_ u2.mem\[181\]\[5\]
+ _01880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_163_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08117_ _03556_ _00022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09097_ _04161_ u2.mem\[22\]\[10\] _04192_ _04195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13455__CLK clknet_leaf_302_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06622__A1 _02044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08048_ _03489_ _03505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09411__I1 u2.mem\[29\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10557__I0 _05101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07178__A2 _02654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10010_ _04764_ _00707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09999_ _04757_ _00703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06386__B1 _01646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06386__C2 _01642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11826__I _05895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06925__A2 _02403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09175__I0 _04164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11961_ _05977_ _01445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06689__A1 u2.mem\[145\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10912_ _05301_ u2.mem\[132\]\[2\] _05319_ _05322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11892_ u2.mem\[192\]\[6\] _03513_ _05937_ _05938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10843_ _05194_ u2.mem\[128\]\[0\] _05278_ _05279_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10378__S _04989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09478__I1 u2.mem\[31\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07638__B1 _03032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13562_ _01441_ clknet_leaf_40_clock u2.mem\[193\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10774_ _05204_ u2.mem\[62\]\[4\] _05237_ _05238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12513_ _00392_ clknet_leaf_162_clock u2.mem\[24\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13493_ _01372_ clknet_leaf_296_clock u2.mem\[185\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12444_ _00323_ clknet_leaf_198_clock u2.mem\[20\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06861__A1 row_select_trans\[0\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08989__I0 _04046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12375_ _00254_ clknet_leaf_59_clock u2.mem\[15\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10905__I _05275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11002__S _05372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10796__I0 _05227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11326_ _05582_ _01205_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06613__A1 _02007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12822__CLK clknet_leaf_83_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11257_ _05540_ _01178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09402__I1 u2.mem\[29\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10548__I0 _05093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07169__A2 _02645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10208_ _04884_ _00785_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11188_ _05495_ _01154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06377__C2 _01653_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10139_ _04844_ _00756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09166__I0 _04151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08913__I0 _04048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11672__S _05801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07877__B1 _02511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12202__CLK clknet_leaf_54_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13328__CLK clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10288__S _04933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06695__A4 _02178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07350_ _02539_ _02825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11276__I1 u2.mem\[154\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06301_ _01798_ _01799_ _01800_ _01805_ _01806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_148_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12352__CLK clknet_leaf_148_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07281_ _02753_ _02754_ _02755_ _02756_ _02757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__13478__CLK clknet_leaf_290_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09020_ _04139_ _04140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06232_ u2.mem\[144\]\[1\] _01671_ _01673_ u2.mem\[182\]\[1\] _01738_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06852__B2 u2.mem\[191\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08780__I mem_address_trans\[4\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06163_ _01638_ _01634_ _01670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_172_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10787__I0 _05218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06094_ _01599_ _01600_ _01601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_100_clock_I clknet_5_11_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09922_ _04712_ u2.mem\[41\]\[13\] _04710_ _04713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10539__I0 _05023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09853_ _04583_ u2.mem\[40\]\[5\] _04666_ _04668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06368__B1 _01683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08804_ _03989_ _04000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_100_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10550__I _04991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09784_ _04617_ _04628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_22_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06996_ _02474_ _02475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09157__I0 _04136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07580__A2 _03049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08735_ _03958_ _00238_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08020__I mem_address_trans\[1\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11582__S _05738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08904__I0 _04039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08666_ _03675_ _03914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08955__I _04094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09321__A3 _03878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09052__S _04155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07617_ _02616_ _03088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08380__I1 u2.mem\[6\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10198__S _04875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08597_ _03870_ _00188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09987__S _04750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07548_ _02414_ _03019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_25_clock_I clknet_5_2_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11267__I1 u2.mem\[154\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10926__S _05327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07479_ u2.mem\[57\]\[6\] _02828_ _02829_ u2.mem\[41\]\[6\] _02952_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09218_ _04251_ _04270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_139_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10490_ _05011_ u2.mem\[55\]\[8\] _05061_ _05062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12845__CLK clknet_leaf_205_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09149_ _04224_ _04122_ _04225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_5_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10725__I _05195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10778__I0 _05209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12160_ _00039_ clknet_leaf_152_clock u2.mem\[2\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11111_ _05448_ _01124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06071__A2 _01565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10661__S _05162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12091_ net23 clknet_2_3__leaf_clock_a inverter_select_trans.A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12995__CLK clknet_leaf_323_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11042_ _05405_ _01098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07020__A1 _02454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12225__CLK clknet_leaf_232_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10950__I0 _05346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09026__I _04144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_302_clock_I clknet_5_16_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12993_ _00872_ clknet_leaf_239_clock u2.mem\[54\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11492__S _05682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08865__I _03709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11944_ _05225_ u2.mem\[193\]\[13\] _05965_ _05967_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10702__I0 _05121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11875_ _03486_ _05926_ _05927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12375__CLK clknet_leaf_59_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10826_ u2.mem\[63\]\[11\] _03525_ _05263_ _05267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11258__I1 u2.mem\[153\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12039__D net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10757_ _03717_ _05227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13545_ _01424_ clknet_leaf_41_clock u2.mem\[192\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07626__A3 _03093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09696__I _04117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13476_ _01355_ clknet_leaf_295_clock u2.mem\[182\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10688_ _05108_ u2.mem\[60\]\[6\] _05179_ _05182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12427_ _00306_ clknet_leaf_178_clock u2.mem\[19\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10769__I0 _05200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12358_ _00237_ clknet_leaf_80_clock u2.mem\[14\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11430__I1 u2.mem\[164\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08105__I _03497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07929__A4 _03393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11309_ _05554_ u2.mem\[156\]\[4\] _05567_ _05573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13000__CLK clknet_leaf_322_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12289_ _00168_ clknet_leaf_165_clock u2.mem\[10\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_343_clock clknet_5_5_0_clock clknet_leaf_343_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_122_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07011__A1 u2.mem\[53\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07165__B _02359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06850_ u2.mem\[185\]\[5\] _02120_ _02122_ u2.mem\[173\]\[5\] _02330_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08976__S _04107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09139__I0 _04167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07562__A2 _03031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06781_ u2.mem\[150\]\[3\] _02047_ _02034_ u2.mem\[174\]\[3\] u2.mem\[181\]\[3\]
+ _02038_ _02263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_110_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08520_ _03824_ u2.mem\[9\]\[11\] _03818_ _03825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12718__CLK clknet_leaf_252_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11497__I1 u2.mem\[168\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_358_clock clknet_5_1_0_clock clknet_leaf_358_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_64_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08451_ _03668_ u2.mem\[8\]\[2\] _03778_ _03781_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07402_ u2.mem\[3\]\[5\] _02801_ _02745_ _02876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08382_ _03727_ _03738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_149_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12868__CLK clknet_leaf_83_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_199_clock_I clknet_5_28_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07333_ u2.mem\[53\]\[4\] _02806_ _02807_ u2.mem\[56\]\[4\] _02808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06825__A1 u2.mem\[171\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06286__C1 _01589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07264_ u2.mem\[27\]\[3\] _02428_ _02436_ u2.mem\[35\]\[3\] _02740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08216__S _03619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09003_ data_in_trans\[1\].data_sync _04126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06215_ _01721_ _01722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10545__I _04986_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07195_ _02572_ _02673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06146_ _01607_ _01629_ _01653_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11421__I1 u2.mem\[163\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_251_clock_I clknet_5_22_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10481__S _05056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06077_ col_select_trans\[2\].data_sync _01584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12248__CLK clknet_leaf_55_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07854__I _02616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09905_ _04682_ _04701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_67_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11185__I0 _05464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09836_ _04657_ _00640_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08886__S _04051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10932__I0 _05307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06979_ _02417_ _02458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_86_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09767_ _04565_ u2.mem\[38\]\[0\] _04618_ _04619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12398__CLK clknet_leaf_179_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08718_ _03917_ u2.mem\[14\]\[5\] _03947_ _03949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09698_ _04121_ _04542_ _04566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_2226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11488__I1 u2.mem\[167\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09550__I0 _04476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08649_ _03725_ _03482_ _03901_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_11660_ _05793_ _01328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07069__A1 _02547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10611_ _05106_ u2.mem\[58\]\[5\] _05136_ _05138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11591_ _05667_ _05750_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_161_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13330_ _01209_ clknet_leaf_3_clock u2.mem\[158\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06933__I _02346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10542_ _05091_ _00912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13261_ _01140_ clknet_leaf_270_clock u2.mem\[147\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10473_ _05052_ _00882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13023__CLK clknet_leaf_249_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12212_ _00091_ clknet_leaf_67_clock u2.mem\[5\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13192_ _01071_ clknet_leaf_276_clock u2.mem\[135\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10376__A1 _04121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12143_ _00022_ clknet_leaf_218_clock u2.mem\[1\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07241__A1 u2.mem\[37\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09369__I0 _04362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13173__CLK clknet_leaf_263_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12074_ data_in_trans\[12\].A clknet_leaf_343_clock data_in_trans\[12\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11025_ _05394_ _05395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_46_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08796__S _03995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06752__B1 _02157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12976_ _00855_ clknet_leaf_249_clock u2.mem\[53\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11927_ _05957_ _01431_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11858_ _05916_ _01403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07004__I _02412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10809_ _05257_ _01013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11100__I0 _05432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11789_ _05873_ _01377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06807__A1 u2.mem\[174\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06807__B2 u2.mem\[181\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13528_ _01407_ clknet_leaf_317_clock u2.mem\[191\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08009__B1 _03462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10365__I _04965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13459_ _01338_ clknet_leaf_345_clock u2.mem\[180\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06000_ u2.driver_mem\[3\] _01508_ _01509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11403__I1 u2.mem\[162\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13516__CLK clknet_leaf_338_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11397__S _05625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_282_clock clknet_5_21_0_clock clknet_leaf_282_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07951_ _01976_ _03246_ _03394_ _03415_ _01491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11196__I _05499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06902_ _02355_ _02380_ _02381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_25_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12540__CLK clknet_leaf_189_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07882_ u2.mem\[14\]\[13\] _02526_ _02528_ u2.mem\[12\]\[13\] _03348_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07535__A2 _02920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06338__A3 _01828_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09621_ _04072_ _04441_ _04521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09780__I0 _04586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06833_ u2.mem\[180\]\[5\] _02042_ _02014_ u2.mem\[172\]\[5\] _02313_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10390__I1 u2.mem\[53\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_297_clock clknet_5_17_0_clock clknet_leaf_297_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09552_ _04147_ _04478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06764_ u2.mem\[194\]\[3\] _02198_ _02199_ u2.mem\[190\]\[3\] _02246_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12690__CLK clknet_5_27_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08503_ _03684_ _03813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09483_ _04384_ u2.mem\[31\]\[12\] _04434_ _04435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06695_ _02172_ _02173_ _02175_ _02178_ _02179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_36_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_220_clock clknet_5_28_0_clock clknet_leaf_220_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08434_ _03710_ u2.mem\[7\]\[12\] _03769_ _03770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08365_ _03657_ u2.mem\[6\]\[0\] _03728_ _03729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13046__CLK clknet_leaf_25_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10476__S _05051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07849__I _02605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07316_ _02781_ _02784_ _02787_ _02790_ _02791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08296_ _03672_ u2.mem\[5\]\[3\] _03660_ _03673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11642__I1 u2.mem\[177\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07066__A4 _02519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_235_clock clknet_5_18_0_clock clknet_leaf_235_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07247_ u2.mem\[28\]\[2\] _02585_ _02587_ u2.mem\[31\]\[2\] _02724_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07471__A1 u2.mem\[14\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07471__B2 u2.mem\[12\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09599__I0 _04478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12070__CLK clknet_leaf_28_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07178_ u2.mem\[44\]\[1\] _02654_ _02655_ u2.mem\[42\]\[1\] _02656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06129_ _01635_ _01636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08271__I0 _03577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11100__S _05434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07584__I _02545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07774__A2 _03091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11158__I0 _05466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09771__I0 _04573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09819_ _04589_ u2.mem\[39\]\[7\] _04644_ _04648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12830_ _00709_ clknet_leaf_220_clock u2.mem\[44\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06928__I _02387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09523__I0 _04384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12761_ _00640_ clknet_leaf_141_clock u2.mem\[39\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11330__I0 _05583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11770__S _05857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11712_ _05824_ _01349_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12692_ _00571_ clknet_leaf_89_clock u2.mem\[35\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11643_ _05782_ _01322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10386__S _04989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06663__I _02147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11574_ _05707_ u2.mem\[173\]\[0\] _05739_ _05740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12413__CLK clknet_leaf_197_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13539__CLK clknet_leaf_34_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07057__A4 _02535_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput17 data_in_a[4] net17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput28 mem_address_a[4] net28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10525_ _05009_ u2.mem\[56\]\[7\] _05078_ _05082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13313_ _01192_ clknet_leaf_349_clock u2.mem\[155\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput39 row_select_a[2] net39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07462__B2 u2.mem\[33\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06804__A4 _02284_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13244_ _01123_ clknet_leaf_291_clock u2.mem\[144\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10456_ _05042_ _00875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11397__I0 _05627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06017__A2 _01517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12563__CLK clknet_leaf_94_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08262__I0 _03568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13175_ _01054_ clknet_leaf_265_clock u2.mem\[132\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10387_ _04996_ _00852_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11010__S _05382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07765__A2 _03072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12126_ _01467_ clknet_leaf_336_clock u2.driver_mem\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_147_clock_I clknet_5_24_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12052__D data_in_trans\[1\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12057_ net17 clknet_2_1__leaf_clock_a data_in_trans\[4\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11008_ _05383_ _01086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09214__I _04150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09514__I0 _04375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08317__I1 u2.mem\[5\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12959_ _00838_ clknet_leaf_155_clock u2.mem\[52\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11321__I0 _05552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13069__CLK clknet_leaf_259_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11680__S _05800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06480_ u2.mem\[0\]\[12\] _01969_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07669__I _02572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12093__CLK clknet_leaf_363_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08150_ _03535_ _03579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11624__I1 u2.mem\[176\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07101_ _02579_ _02580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07453__A1 _02905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06256__A2 _01715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08081_ _03528_ _03529_ _03530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12906__CLK clknet_leaf_141_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07032_ _02510_ _02511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08253__I0 _03559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07756__A2 _03213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08983_ _04111_ _00333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07934_ _03395_ _03396_ _03397_ _03398_ _03399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_29_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09325__S _04336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07865_ _01969_ _03246_ _03286_ _03331_ _01489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11560__I0 _05707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09604_ _04482_ u2.mem\[34\]\[8\] _04511_ _04512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06816_ u2.mem\[153\]\[4\] _02196_ _02200_ u2.mem\[160\]\[4\] _02297_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07796_ u2.mem\[1\]\[12\] _03261_ _03262_ u2.mem\[7\]\[12\] _03263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09505__I0 _04366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_349_clock_I clknet_5_4_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09535_ _04466_ _00530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06747_ _02227_ _02228_ _02229_ _02230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_43_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10115__I1 u2.mem\[46\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09466_ _04425_ _00502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06678_ _02049_ _02074_ _02113_ _02162_ _02163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__11863__I1 u2.mem\[191\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07141__B1 _02619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08417_ _03760_ _00118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09397_ _04163_ _04382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07579__I _02516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_174_clock clknet_5_27_0_clock clknet_leaf_174_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08348_ _03714_ _03715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12586__CLK clknet_leaf_115_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07444__B2 u2.mem\[19\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08279_ _03658_ _03544_ _03633_ _03659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_10310_ _04895_ u2.mem\[51\]\[4\] _04949_ _04950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11290_ _05550_ u2.mem\[155\]\[2\] _05559_ _05562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11379__I0 _05583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_189_clock clknet_5_31_0_clock clknet_leaf_189_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_152_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10241_ _04907_ u2.mem\[49\]\[9\] _04905_ _04908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08244__I0 _03550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10051__I0 _04788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07747__A2 _03114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10172_ _03983_ _04863_ _04864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_79_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_112_clock clknet_5_14_0_clock clknet_leaf_112_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_121_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11551__I0 _05715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13211__CLK clknet_leaf_287_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06183__A1 u2.mem\[170\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09034__I _04150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06183__B2 u2.mem\[156\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_127_clock clknet_5_15_0_clock clknet_leaf_127_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_28_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12813_ _00692_ clknet_leaf_201_clock u2.mem\[43\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11303__I0 _05548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12744_ _00623_ clknet_leaf_50_clock u2.mem\[38\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11854__I1 u2.mem\[190\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13361__CLK clknet_leaf_355_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06486__A2 _01933_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12675_ _00554_ clknet_leaf_86_clock u2.mem\[34\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_73_clock_I clknet_5_8_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12929__CLK clknet_leaf_233_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11626_ _05750_ u2.mem\[176\]\[1\] _05771_ _05773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_1553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06238__A2 _01676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07435__B2 u2.mem\[11\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11557_ _05605_ _05729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_156_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10508_ _04224_ _05071_ _05072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_170_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11488_ _05674_ u2.mem\[167\]\[3\] _05683_ _05687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10990__A1 _04249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09188__A1 _03901_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13227_ _01106_ clknet_leaf_279_clock u2.mem\[141\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10439_ _04995_ u2.mem\[54\]\[2\] _05030_ _05033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07199__B1 _02582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07738__A2 _03021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_298_clock_I clknet_5_17_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13158_ _01037_ clknet_leaf_269_clock u2.mem\[129\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12309__CLK clknet_leaf_100_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10593__I1 u2.mem\[57\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12109_ _01492_ clknet_leaf_140_clock u2.active_mem\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13089_ _00968_ clknet_leaf_241_clock u2.mem\[60\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09145__S _04218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10345__I1 u2.mem\[52\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07650_ _02520_ _03120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12459__CLK clknet_leaf_179_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_350_clock_I clknet_5_4_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06601_ _02023_ _02033_ _02086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07581_ _03046_ _03047_ _03048_ _03051_ _03052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_80_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09320_ _04332_ _00449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09879__I _04682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06532_ _02016_ _01986_ _02017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11845__I1 u2.mem\[190\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_91_clock clknet_5_10_0_clock clknet_leaf_91_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09251_ _04256_ u2.mem\[26\]\[2\] _04290_ _04293_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06463_ u2.mem\[192\]\[8\] _01931_ _01956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07674__B2 u2.mem\[31\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08202_ _03550_ u2.mem\[3\]\[2\] _03609_ _03612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09182_ _04174_ u2.mem\[24\]\[14\] _04241_ _04244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06394_ _01888_ _01889_ _01890_ _01895_ _01896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_159_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08133_ _03567_ _00027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08474__I0 _03710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08064_ _03489_ _03517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07015_ _02413_ _02491_ _02492_ _02493_ _02494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_31_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10553__I _04994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07729__A2 _03088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06401__A2 _01719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08966_ _04096_ _04102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_input31_I mem_address_a[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07917_ u2.mem\[3\]\[14\] _03267_ _03211_ _03382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08897_ _04050_ _04061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_116_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_44_clock clknet_5_6_0_clock clknet_leaf_44_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_56_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07848_ u2.mem\[52\]\[12\] _03313_ _03314_ u2.mem\[21\]\[12\] _03315_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06165__A1 _01665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13384__CLK clknet_leaf_301_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07779_ _02360_ _03246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09518_ _04380_ u2.mem\[32\]\[10\] _04453_ _04456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08693__I _03905_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_59_clock clknet_5_12_0_clock clknet_leaf_59_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_10790_ _05246_ _01005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09449_ _04414_ _00496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10728__I _05004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_12460_ _00339_ clknet_leaf_196_clock u2.mem\[21\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11411_ _04071_ _05606_ _05637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_123_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12391_ _00270_ clknet_leaf_134_clock u2.mem\[16\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08465__I0 _03693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07968__A2 _02526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11342_ _05593_ u2.mem\[158\]\[4\] _05584_ _05594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06941__I _02419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08090__A1 _03535_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11559__I _05730_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11273_ _05550_ u2.mem\[154\]\[2\] _05546_ _05551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09029__I data_in_trans\[6\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08917__A1 _04072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10224_ _04886_ _04896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09965__I0 _04716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13012_ _00891_ clknet_leaf_31_clock u2.mem\[55\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11772__I0 _05835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10155_ _04853_ _00763_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09717__I0 _04579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12601__CLK clknet_leaf_116_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10086_ _04608_ _04813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06156__A1 _01617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09699__I _04566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11827__I1 u2.mem\[189\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10988_ _05352_ u2.mem\[136\]\[5\] _05364_ _05371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12727_ _00606_ clknet_leaf_43_clock u2.mem\[37\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06459__A2 _01942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08108__I _03500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12658_ _00537_ clknet_leaf_224_clock u2.mem\[33\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13107__CLK clknet_leaf_20_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07012__I _02430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08456__I0 _03676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10574__S _05113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11609_ _05762_ _01308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12589_ _00468_ clknet_leaf_187_clock u2.mem\[29\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08081__A1 _03528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12131__CLK clknet_leaf_35_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13257__CLK clknet_leaf_312_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09956__I0 _04707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07187__A3 _02653_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08820_ _03939_ u2.mem\[16\]\[15\] _04005_ _04009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06395__A1 u2.mem\[190\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06395__B2 u2.mem\[194\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12281__CLK clknet_leaf_119_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09708__I0 _04573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08751_ _03967_ _00245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11515__I0 _05671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07702_ u2.mem\[50\]\[10\] _03111_ _03112_ u2.mem\[51\]\[10\] _03171_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08682_ _03925_ _00218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07633_ u2.mem\[40\]\[9\] _03018_ _03019_ u2.mem\[30\]\[9\] _03103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07895__B2 u2.mem\[31\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11932__I _05949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07564_ u2.mem\[3\]\[8\] _03034_ _02978_ _03035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11999__CLK clknet_leaf_28_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09303_ _04312_ _04323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06515_ _01999_ _02000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07495_ _02964_ _02965_ _02966_ _02967_ _02968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09234_ _04170_ _04281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06446_ _01927_ _01942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09165_ _04234_ _00392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08447__I0 _03657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06377_ u2.mem\[189\]\[5\] _01650_ _01652_ u2.mem\[176\]\[5\] u2.mem\[172\]\[5\]
+ _01653_ _01879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_33_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10254__I0 _04916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08116_ _03554_ u2.mem\[1\]\[4\] _03555_ _03556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07857__I _02611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09096_ _04194_ _00363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08611__A3 _03878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06083__B1 _01589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08047_ _01809_ _03490_ _03504_ _00004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06622__A2 _02104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09947__I0 _04698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12624__CLK clknet_leaf_168_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11754__I0 _05831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_21_clock_I clknet_5_2_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09998_ _04712_ u2.mem\[43\]\[13\] _04755_ _04757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06386__B2 u2.mem\[165\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07583__B1 _02900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06925__A3 _02383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08949_ _04091_ _00319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09175__I1 u2.mem\[24\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06138__A1 _01570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11960_ _05911_ u2.mem\[194\]\[3\] _05975_ _05977_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10911_ _05321_ _01051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06001__I _01502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07886__A1 _03336_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10659__S _05162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11891_ _05928_ _05937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06936__I _02414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10842_ _05277_ _05278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_leaf_246_clock_I clknet_5_22_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12004__CLK clknet_leaf_40_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08129__S _03564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09312__I _04312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13561_ _01440_ clknet_leaf_32_clock u2.mem\[193\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10773_ _05231_ _05237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_164_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12512_ _00391_ clknet_leaf_162_clock u2.mem\[24\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13492_ _01371_ clknet_leaf_292_clock u2.mem\[185\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12154__CLK clknet_leaf_56_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12443_ _00322_ clknet_leaf_199_clock u2.mem\[20\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08438__I0 _03719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08989__I1 u2.mem\[20\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06671__I _02155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08063__A1 _01951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12374_ _00253_ clknet_leaf_78_clock u2.mem\[15\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10796__I1 u2.mem\[62\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11325_ _05556_ u2.mem\[157\]\[5\] _05575_ _05582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06613__A2 _02080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09938__I0 _04689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11256_ _05508_ u2.mem\[153\]\[2\] _05537_ _05540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11745__I0 _05837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10207_ _04817_ u2.mem\[48\]\[15\] _04880_ _04884_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10921__I _05326_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11187_ _05466_ u2.mem\[149\]\[2\] _05492_ _05495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06377__A1 u2.mem\[189\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10138_ _04788_ u2.mem\[47\]\[2\] _04841_ _04844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11953__S _05972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12060__D data_in_trans\[5\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10069_ _04591_ _04801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07007__I _02485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09423__S _04396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08913__I1 u2.mem\[18\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08677__I0 _03921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06300_ u2.mem\[147\]\[2\] _01676_ _01680_ u2.mem\[169\]\[2\] _01804_ _01805_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_91_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07280_ u2.mem\[43\]\[3\] _02515_ _02517_ u2.mem\[20\]\[3\] _02756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06301__A1 _01798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06231_ u2.mem\[158\]\[1\] _01728_ _01729_ u2.mem\[151\]\[1\] _01736_ _01737_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08429__I0 _03702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06852__A2 _02150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07677__I _02597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06581__I _02065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06162_ _01655_ _01662_ _01668_ _01669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12647__CLK clknet_leaf_114_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10936__A1 _04180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11984__I0 _05227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07801__A1 u2.mem\[3\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06093_ _01587_ _01600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09892__I _04682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09921_ _04608_ _04712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12797__CLK clknet_leaf_220_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08601__I0 _03826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09852_ _04667_ _00646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_195_clock_I clknet_5_31_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06368__A1 u2.mem\[191\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06368__B2 u2.mem\[179\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08803_ _03999_ _00265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08301__I _03659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09783_ _04627_ _00617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_06995_ _02388_ _02390_ _02384_ _02473_ _02474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08734_ _03932_ u2.mem\[14\]\[12\] _03957_ _03958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12027__CLK clknet_2_0__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08665_ _03913_ _00213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07868__B2 u2.mem\[30\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07616_ u2.mem\[5\]\[8\] _02920_ _02921_ u2.mem\[38\]\[8\] _03087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08596_ _03822_ u2.mem\[11\]\[10\] _03867_ _03870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12177__CLK clknet_leaf_218_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07547_ _02405_ _03018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08668__I0 _03914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07478_ u2.mem\[37\]\[6\] _02825_ _02826_ u2.mem\[59\]\[6\] _02951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09217_ _04153_ _04269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06429_ _01918_ _01929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07587__I _02539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09093__I0 _04154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09148_ _04223_ _04224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_108_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13572__CLK clknet_leaf_20_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09079_ _04132_ u2.mem\[22\]\[2\] _04182_ _04185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10942__S _05337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11110_ _05426_ u2.mem\[144\]\[2\] _05445_ _05448_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12090_ output_active_trans.A clknet_leaf_303_clock output_active_trans.data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11041_ _05380_ u2.mem\[140\]\[0\] _05404_ _05405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10741__I _03696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11104__A1 _03487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12992_ _00871_ clknet_leaf_240_clock u2.mem\[54\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11943_ _05966_ _01438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07859__B2 u2.mem\[4\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06666__I _02150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11874_ _03477_ mem_address_trans\[5\].data_sync _05925_ _05926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_2975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09042__I data_in_trans\[9\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10825_ _05266_ _01020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09977__I _04739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10466__I0 _05025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13544_ _01423_ clknet_leaf_32_clock u2.mem\[192\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10756_ _05226_ _00991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06834__A2 _02311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13475_ _01354_ clknet_leaf_295_clock u2.mem\[182\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10687_ _05181_ _00967_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10218__I0 _04891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11013__S _05382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12426_ _00305_ clknet_leaf_112_clock u2.mem\[18\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09084__I0 _04140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11948__S _05965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12055__D net16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08831__I0 _04017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12357_ _00236_ clknet_leaf_80_clock u2.mem\[14\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06598__A1 u2.mem\[165\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06598__B2 u2.mem\[163\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11308_ _05572_ _01197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12288_ _00167_ clknet_leaf_165_clock u2.mem\[10\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11747__I _05768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11239_ _05530_ _01170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09217__I _04153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08121__I _03513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07011__A2 _02486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06780_ u2.mem\[155\]\[3\] _02029_ _02262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06770__A1 u2.mem\[167\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09153__S _04226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06770__B2 u2.mem\[183\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08898__I0 _04032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13445__CLK clknet_leaf_350_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08450_ _03780_ _00131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07401_ u2.mem\[16\]\[5\] _02798_ _02799_ u2.mem\[33\]\[5\] _02875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08381_ _03737_ _00105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10457__I0 _05016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07332_ _02488_ _02807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07078__A2 _02554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06286__B1 _01572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07263_ u2.mem\[40\]\[3\] _02406_ _02415_ u2.mem\[30\]\[3\] _02739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09002_ _04125_ _00338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06214_ _01678_ _01582_ _01613_ _01721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__08027__A1 _03480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09075__I0 _04119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07194_ _02668_ _02669_ _02670_ _02671_ _02672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_69_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06145_ _01651_ _01652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07250__A2 _02591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06076_ _01582_ _01576_ _01583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_160_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11709__I0 _05796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09904_ _04591_ _04700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11185__I1 u2.mem\[149\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07002__A2 _02480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09835_ _04612_ u2.mem\[39\]\[14\] _04654_ _04657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08031__I _03491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08966__I _04096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09766_ _04617_ _04618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_73_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06978_ _02456_ _02457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08717_ _03948_ _00230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08889__I0 _04023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09697_ _04564_ _04565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09998__S _04755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10002__S _04755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08648_ _03656_ _03900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06513__A1 row_select_trans\[5\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07710__B1 _03050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12812__CLK clknet_leaf_201_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08579_ _03860_ _00180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10448__I0 _05007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_10610_ _05137_ _00934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07069__A2 _02371_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11590_ _05749_ _01302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06277__B1 _01658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06277__C2 u2.mem\[181\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10541_ _05025_ u2.mem\[56\]\[14\] _05088_ _05091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08206__I _03608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13260_ _01139_ clknet_leaf_295_clock u2.mem\[146\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10472_ _04987_ u2.mem\[55\]\[0\] _05051_ _05052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11948__I0 _05229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12211_ _00090_ clknet_leaf_65_clock u2.mem\[5\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11768__S _05857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13191_ _01070_ clknet_leaf_279_clock u2.mem\[135\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10376__A2 _04964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10620__I0 _05115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12142_ _00021_ clknet_leaf_211_clock u2.mem\[1\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13318__CLK clknet_leaf_301_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07241__A2 _02540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_0_clock_a clock_a clknet_0_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_2_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09369__I1 u2.mem\[29\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10471__I _05050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12073_ net10 clknet_2_1__leaf_clock_a data_in_trans\[12\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09037__I data_in_trans\[8\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11024_ _04311_ _05363_ _05394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_89_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12342__CLK clknet_leaf_78_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13468__CLK clknet_leaf_346_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06752__A1 u2.mem\[146\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12975_ _00854_ clknet_leaf_249_clock u2.mem\[53\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11926_ _05915_ u2.mem\[193\]\[5\] _05955_ _05957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12492__CLK clknet_leaf_190_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11857_ _05915_ u2.mem\[190\]\[5\] _05904_ _05916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10847__S _05278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_143_clock_I clknet_5_24_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10439__I0 _04995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10808_ u2.mem\[63\]\[3\] _03503_ _05253_ _05257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08317__S _03677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11788_ _05872_ u2.mem\[186\]\[3\] _05866_ _05873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13527_ _01406_ clknet_leaf_316_clock u2.mem\[191\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10739_ _05213_ u2.mem\[61\]\[8\] _05214_ _05215_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08009__A1 u2.active_mem\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09057__I0 _04167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08009__B2 u2.active_mem\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13458_ _01337_ clknet_leaf_306_clock u2.mem\[179\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07480__A2 _02950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11939__I0 _05220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11678__S _05801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12409_ _00288_ clknet_leaf_122_clock u2.mem\[17\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13389_ _01268_ clknet_leaf_355_clock u2.mem\[168\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07768__B1 _03078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10611__I0 _05106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10381__I _04991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07950_ _03399_ _03404_ _03409_ _03414_ _03415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_155_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06991__A1 _02466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06901_ _02352_ _02341_ _02342_ _02379_ _02380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA_clkbuf_leaf_68_clock_I clknet_5_9_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07881_ u2.mem\[44\]\[13\] _02521_ _02523_ u2.mem\[42\]\[13\] _03347_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09620_ _04520_ _00561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06338__A4 _01841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08786__I _03989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06832_ u2.mem\[176\]\[5\] _02004_ _02020_ u2.mem\[189\]\[5\] _02312_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07940__B1 _02598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09551_ _04477_ _00535_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06763_ u2.mem\[154\]\[3\] _02225_ _02226_ u2.mem\[162\]\[3\] _02245_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08502_ _03812_ _00151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09482_ _04418_ _04434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07299__A2 _02617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06694_ u2.mem\[149\]\[1\] _02176_ _02177_ u2.mem\[175\]\[1\] _02178_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08433_ _03753_ _03769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_52_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12985__CLK clknet_leaf_319_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08364_ _03727_ _03728_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_51_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09410__I _04176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07315_ u2.mem\[27\]\[4\] _02788_ _02789_ u2.mem\[35\]\[4\] _02790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10556__I _04997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08295_ _03671_ _03672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07246_ u2.mem\[9\]\[2\] _02580_ _02582_ u2.mem\[25\]\[2\] _02723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09048__I0 _04161_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12215__CLK clknet_leaf_53_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07471__A2 _02890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07177_ _02522_ _02655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10492__S _05061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_345_clock_I clknet_5_5_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06128_ _01552_ _01634_ _01635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10602__I0 _05097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07223__A2 _02457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08271__I1 u2.mem\[4\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12365__CLK clknet_leaf_210_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06059_ _01556_ _01566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11158__I1 u2.mem\[147\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09818_ _04647_ _00632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08696__I _03714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09771__I1 u2.mem\[38\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06734__A1 u2.mem\[159\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06734__B2 u2.mem\[149\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09749_ _04604_ _04605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09523__I1 u2.mem\[32\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12760_ _00639_ clknet_leaf_51_clock u2.mem\[39\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11330__I1 u2.mem\[158\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11711_ _05798_ u2.mem\[181\]\[5\] _05817_ _05824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06498__B1 _01970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12691_ _00570_ clknet_leaf_89_clock u2.mem\[35\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11850__I _03670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11642_ _05752_ u2.mem\[177\]\[2\] _05779_ _05782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11094__I0 _05426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_342_clock clknet_5_5_0_clock clknet_leaf_342_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11573_ _05738_ _05739_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_52_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput18 data_in_a[5] net18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13312_ _01191_ clknet_leaf_348_clock u2.mem\[155\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10524_ _05081_ _00904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput29 mem_address_a[5] net29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13140__CLK clknet_leaf_22_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13243_ _01122_ clknet_leaf_291_clock u2.mem\[144\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12708__CLK clknet_leaf_68_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10455_ _05014_ u2.mem\[54\]\[9\] _05040_ _05042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11397__I1 u2.mem\[162\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_357_clock clknet_5_1_0_clock clknet_leaf_357_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_151_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07214__A2 _02622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13174_ _01053_ clknet_leaf_275_clock u2.mem\[132\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08262__I1 u2.mem\[4\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10386_ _04995_ u2.mem\[53\]\[2\] _04989_ _04996_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12125_ _01466_ clknet_leaf_334_clock u2.driver_mem\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13290__CLK clknet_leaf_354_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12858__CLK clknet_leaf_129_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12056_ data_in_trans\[3\].A clknet_leaf_288_clock data_in_trans\[3\].data_sync vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11007_ _05380_ u2.mem\[138\]\[0\] _05382_ _05383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06725__A1 u2.mem\[184\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09514__I1 u2.mem\[32\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12958_ _00837_ clknet_leaf_197_clock u2.mem\[52\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11321__I1 u2.mem\[157\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11909_ u2.mem\[192\]\[14\] _03533_ _05928_ _05947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10577__S _05113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12889_ _00768_ clknet_leaf_51_clock u2.mem\[47\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_294_clock_I clknet_5_20_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09278__I0 _04283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12238__CLK clknet_leaf_211_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09230__I _04166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07100_ _02577_ _02578_ _02552_ _02455_ _02579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_105_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08080_ _03493_ _03529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07453__A2 _02912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07031_ _02487_ _02496_ _02497_ _02468_ _02510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_174_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07205__A2 _02591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09450__I0 _04391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07756__A3 _03218_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08982_ _04039_ u2.mem\[20\]\[11\] _04107_ _04111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06964__A1 _02398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09606__S _04511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09202__I0 _04258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07933_ u2.mem\[57\]\[14\] _03294_ _03295_ u2.mem\[41\]\[14\] _03398_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08705__A2 _03726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07864_ _03297_ _03308_ _03319_ _03330_ _03331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_83_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09603_ _04500_ _04511_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_99_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11560__I1 u2.mem\[172\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06815_ u2.mem\[194\]\[4\] _02198_ _02199_ u2.mem\[190\]\[4\] _02296_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07795_ _02470_ _03262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09505__I1 u2.mem\[32\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09534_ _04463_ u2.mem\[33\]\[0\] _04465_ _04466_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06746_ u2.mem\[148\]\[2\] _02128_ _02130_ u2.mem\[152\]\[2\] _02229_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09465_ _04366_ u2.mem\[31\]\[4\] _04424_ _04425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10487__S _05056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06677_ _02118_ _02124_ _02140_ _02161_ _02162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_24_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08416_ _03676_ u2.mem\[7\]\[4\] _03759_ _03760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09269__I0 _04274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09396_ _04381_ _00476_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07692__A2 _03099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13163__CLK clknet_leaf_274_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08347_ _03713_ _03714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08278_ _03541_ _03658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_138_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07229_ u2.mem\[54\]\[2\] _02648_ _02649_ u2.mem\[55\]\[2\] _02706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07595__I _02564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11379__I1 u2.mem\[161\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10240_ _04595_ _04907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09441__I0 _04382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06404__B1 _01693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10171_ _04862_ _04863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10950__S _05337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06955__A1 _02401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09516__S _04453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06004__I _01512_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11000__I0 _05349_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06939__I _02417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06707__A1 u2.mem\[155\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06707__B2 u2.mem\[174\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11551__I1 u2.mem\[171\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12812_ _00691_ clknet_leaf_201_clock u2.mem\[43\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09251__S _04290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11303__I1 u2.mem\[156\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13506__CLK clknet_leaf_330_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12743_ _00622_ clknet_leaf_53_clock u2.mem\[38\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08180__I0 _03568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12674_ _00553_ clknet_leaf_154_clock u2.mem\[34\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_281_clock clknet_5_21_0_clock clknet_leaf_281_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_16_clock_I clknet_5_2_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09050__I data_in_trans\[11\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11625_ _05772_ _01314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12530__CLK clknet_leaf_166_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11556_ _05728_ _01289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10507_ _04862_ _05071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06789__A4 _02270_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_296_clock clknet_5_17_0_clock clknet_leaf_296_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11487_ _05686_ _01262_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05997__A2 row_col_select_trans.data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13226_ _01105_ clknet_leaf_279_clock u2.mem\[141\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09432__I0 _04373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12680__CLK clknet_leaf_129_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10438_ _05032_ _00867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12063__D net20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13157_ _01036_ clknet_leaf_269_clock u2.mem\[129\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10860__S _05287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10369_ _04983_ _00847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12108_ _01491_ clknet_leaf_135_clock u2.active_mem\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13088_ _00967_ clknet_leaf_245_clock u2.mem\[60\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12039_ net2 clknet_2_2__leaf_clock_a col_select_trans\[1\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_234_clock clknet_5_18_0_clock clknet_leaf_234_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06174__A2 _01599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06600_ _02084_ _02085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07580_ u2.mem\[43\]\[8\] _03049_ _03050_ u2.mem\[20\]\[8\] _03051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_19_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12060__CLK clknet_leaf_300_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13186__CLK clknet_leaf_276_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06531_ _01984_ _02016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_94_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08171__I0 _03559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09250_ _04292_ _00419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_249_clock clknet_5_22_0_clock clknet_leaf_249_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_21_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06462_ _01914_ _01955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07674__A2 _03072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08201_ _03611_ _00051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11058__I0 _05384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09181_ _04243_ _00399_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06393_ u2.mem\[166\]\[5\] _01592_ _01597_ u2.mem\[161\]\[5\] _01894_ _01895_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_18_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09895__I _04582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08132_ _03566_ u2.mem\[1\]\[9\] _03564_ _03567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08063_ _01951_ _03505_ _03516_ _00008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07977__A3 _03439_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07014_ _02401_ _02403_ _02392_ _02493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_108_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08304__I _03510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09423__I0 _04364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08965_ _04101_ _00325_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08240__S _03635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07916_ u2.mem\[16\]\[14\] _03264_ _03265_ u2.mem\[33\]\[14\] _03381_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08896_ _04060_ _00297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12403__CLK clknet_leaf_108_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input24_I mem_address_a[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13529__CLK clknet_leaf_316_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07847_ _02602_ _03314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06165__A2 _01591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07778_ _01966_ _03013_ _03224_ _03245_ _01488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09517_ _04455_ _00523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06729_ u2.mem\[176\]\[2\] _02004_ _02020_ u2.mem\[189\]\[2\] _02212_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12553__CLK clknet_leaf_119_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08162__I0 _03550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11106__S _05445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_09448_ _04389_ u2.mem\[30\]\[14\] _04411_ _04414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07665__A2 _03055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09379_ _04369_ u2.mem\[29\]\[5\] _04367_ _04370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11410_ _05636_ _01235_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12390_ _00269_ clknet_leaf_77_clock u2.mem\[16\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08465__I1 u2.mem\[8\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11341_ _05513_ _05593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10744__I _03700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11272_ _05507_ _05550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_1424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_242_clock_I clknet_5_19_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13059__CLK clknet_leaf_27_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13011_ _00890_ clknet_leaf_323_clock u2.mem\[55\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10223_ _04578_ _04895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11772__I1 u2.mem\[185\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07050__B1 _02528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10154_ _04804_ u2.mem\[47\]\[9\] _04851_ _04853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10085_ _04812_ _00734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12083__CLK clknet_leaf_363_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06156__A2 _01619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11288__I0 _05548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10987_ _05370_ _01078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11016__S _05382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12726_ _00605_ clknet_leaf_72_clock u2.mem\[37\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12058__D data_in_trans\[4\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12657_ _00536_ clknet_leaf_224_clock u2.mem\[33\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11608_ _05746_ u2.mem\[175\]\[0\] _05761_ _05762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12588_ _00467_ clknet_leaf_190_clock u2.mem\[29\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08456__I1 u2.mem\[8\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11539_ _05718_ _01282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10654__I _05151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09405__I0 _04387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08124__I _03515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13209_ _01088_ clknet_leaf_281_clock u2.mem\[138\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11912__A1 _01981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12426__CLK clknet_leaf_112_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07187__A4 _02664_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06395__A2 _01702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08750_ _03912_ u2.mem\[15\]\[3\] _03963_ _03967_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09708__I1 u2.mem\[37\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_173_clock clknet_5_27_0_clock clknet_leaf_173_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_97_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11515__I1 u2.mem\[169\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07701_ _03166_ _03167_ _03168_ _03169_ _03170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_6_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08681_ _03923_ u2.mem\[13\]\[8\] _03924_ _03925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08392__I0 _03710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07632_ u2.mem\[32\]\[9\] _03015_ _03016_ u2.mem\[2\]\[9\] _03102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11279__I0 _05554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_188_clock clknet_5_31_0_clock clknet_leaf_188_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07563_ _02479_ _03034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09302_ _04322_ _00441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06514_ _01998_ _01999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07494_ u2.mem\[6\]\[6\] _02861_ _02862_ u2.mem\[47\]\[6\] _02967_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07647__A2 _03039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07203__I _02597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_191_clock_I clknet_5_31_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09233_ _04280_ _00414_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06855__B1 _02143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06445_ u2.mem\[192\]\[5\] _01931_ _01941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10765__S _05232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_111_clock clknet_5_14_0_clock clknet_leaf_111_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_21_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09164_ _04148_ u2.mem\[24\]\[6\] _04231_ _04234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06376_ _01877_ _01878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08115_ _03545_ _03555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_135_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09095_ _04158_ u2.mem\[22\]\[9\] _04192_ _04194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06083__A1 u2.mem\[177\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07280__B1 _02517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06083__B2 u2.mem\[168\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08046_ _03503_ _03494_ _03504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_126_clock clknet_5_15_0_clock clknet_leaf_126_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_134_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11754__I1 u2.mem\[184\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13351__CLK clknet_leaf_361_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09997_ _04756_ _00702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08948_ _04044_ u2.mem\[19\]\[13\] _04089_ _04091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12919__CLK clknet_leaf_125_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08879_ _04050_ _04051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_3825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08383__I0 _03693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10910_ _05299_ u2.mem\[132\]\[1\] _05319_ _05321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07886__A2 _03341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11890_ _05936_ _01415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10841_ _03983_ _05276_ _05277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_71_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08135__I0 _03568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13560_ _01439_ clknet_leaf_32_clock u2.mem\[193\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07638__A2 _03031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10772_ _05236_ _00997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09883__I0 _04685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12511_ _00390_ clknet_leaf_162_clock u2.mem\[24\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06846__B1 _02137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13491_ _01370_ clknet_leaf_292_clock u2.mem\[185\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10675__S _05174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06310__A2 _01811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12442_ _00321_ clknet_leaf_128_clock u2.mem\[19\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06952__I _02430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11442__I0 _05623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12373_ _00252_ clknet_leaf_79_clock u2.mem\[15\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12449__CLK clknet_leaf_159_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11324_ _05581_ _01204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11255_ _05539_ _01177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08879__I _04050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11745__I1 u2.mem\[183\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10206_ _04883_ _00784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_90_clock clknet_5_8_0_clock clknet_leaf_90_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11186_ _05494_ _01153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07574__A1 _03037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12599__CLK clknet_leaf_113_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10137_ _04843_ _00755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09704__S _04567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10068_ _04800_ _00729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08374__I0 _03676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07877__A2 _02509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12709_ _00588_ clknet_leaf_27_clock u2.mem\[36\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13224__CLK clknet_leaf_286_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06301__A2 _01799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06230_ _01730_ _01733_ _01735_ _01736_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_31_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_43_clock clknet_5_6_0_clock clknet_leaf_43_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10384__I _04130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06161_ u2.mem\[180\]\[0\] _01664_ _01667_ u2.mem\[150\]\[0\] _01668_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_157_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06092_ _01546_ _01560_ _01599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_117_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13374__CLK clknet_leaf_355_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09920_ _04711_ _00670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_58_clock clknet_5_12_0_clock clknet_leaf_58_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_98_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09851_ _04579_ u2.mem\[40\]\[4\] _04666_ _04667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_138_clock_I clknet_5_13_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06368__A2 _01681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08802_ _03921_ u2.mem\[16\]\[7\] _03995_ _03999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09782_ _04589_ u2.mem\[38\]\[7\] _04623_ _04627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_06994_ _02412_ _02473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_86_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08733_ _03941_ _03957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_38_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08365__I0 _03657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08664_ _03912_ u2.mem\[13\]\[3\] _03906_ _03913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07615_ _03076_ _03079_ _03082_ _03085_ _03086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_1708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10872__A1 _05295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10559__I _05000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08595_ _03869_ _00187_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07546_ u2.mem\[32\]\[8\] _03015_ _03016_ u2.mem\[2\]\[8\] _03017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08029__I _03489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11672__I0 _05786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07477_ u2.mem\[60\]\[6\] _02822_ _02823_ u2.mem\[62\]\[6\] _02950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09216_ _04268_ _00409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06428_ _01927_ _01928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09617__I0 _04496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09147_ _03629_ _03749_ _03775_ _04223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_147_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06359_ _01854_ _01855_ _01856_ _01861_ _01862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_30_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09078_ _04184_ _00355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08029_ _03489_ _03490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08699__I _03718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12741__CLK clknet_leaf_70_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11040_ _05403_ _05404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_39_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07108__I _02586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12991_ _00870_ clknet_leaf_239_clock u2.mem\[54\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11853__I _03674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11104__A2 _05443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11942_ _05222_ u2.mem\[193\]\[12\] _05965_ _05966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10163__I0 _04813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06947__I _02412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11873_ mem_address_trans\[6\].data_sync mem_address_trans\[7\].data_sync _05925_
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13247__CLK clknet_leaf_272_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12121__CLK clknet_leaf_328_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10824_ u2.mem\[63\]\[10\] _03523_ _05263_ _05266_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13543_ _01422_ clknet_leaf_32_clock u2.mem\[192\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10755_ _05225_ u2.mem\[61\]\[13\] _05223_ _05226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12271__CLK clknet_leaf_166_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09608__I0 _04487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06295__B2 u2.mem\[185\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13474_ _01353_ clknet_leaf_293_clock u2.mem\[182\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13397__CLK clknet_leaf_307_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10686_ _05106_ u2.mem\[60\]\[5\] _05179_ _05181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12425_ _00304_ clknet_leaf_128_clock u2.mem\[18\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11415__I0 _05627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07244__B1 _02674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12356_ _00235_ clknet_leaf_80_clock u2.mem\[14\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08603__S _03872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11307_ _05552_ u2.mem\[156\]\[3\] _05568_ _05572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12287_ _00166_ clknet_leaf_164_clock u2.mem\[10\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11989__CLK clknet_leaf_318_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11238_ _05500_ u2.mem\[152\]\[0\] _05529_ _05530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11964__S _05975_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12071__D net9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11169_ _05460_ u2.mem\[148\]\[0\] _05484_ _05485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07018__I _02432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10154__I0 _04804_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07400_ u2.mem\[1\]\[5\] _02795_ _02796_ u2.mem\[7\]\[5\] _02874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08380_ _03689_ u2.mem\[6\]\[7\] _03733_ _03737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07331_ _02485_ _02806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_64_clock_I clknet_5_9_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06286__A1 u2.mem\[158\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07262_ u2.mem\[32\]\[3\] _02386_ _02396_ u2.mem\[2\]\[3\] _02738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_91_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06286__B2 u2.mem\[151\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09001_ _04119_ u2.mem\[21\]\[0\] _04124_ _04125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11406__I0 _05633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06213_ _01719_ _01720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08027__A2 _03487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07193_ u2.mem\[57\]\[1\] _02554_ _02556_ u2.mem\[41\]\[1\] _02671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12764__CLK clknet_leaf_203_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07235__B1 _02661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06144_ _01582_ _01634_ _01651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_156_1506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06589__A2 _02063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07786__B2 u2.mem\[30\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10842__I _05277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06075_ _01581_ _01582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11709__I1 u2.mem\[181\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_289_clock_I clknet_5_20_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09903_ _04699_ _00665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06033__S _01541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07538__A1 u2.mem\[6\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09834_ _04656_ _00639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09765_ _04180_ _04542_ _04617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06977_ _02451_ _02452_ _02453_ _02455_ _02456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__12144__CLK clknet_leaf_226_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08338__I0 _03706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06761__A2 _02241_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08716_ _03914_ u2.mem\[14\]\[4\] _03947_ _03948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09696_ _04117_ _04564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10145__I0 _04795_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_341_clock_I clknet_5_5_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08647_ _03899_ _00209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07710__B2 u2.mem\[20\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12294__CLK clknet_leaf_101_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08578_ _03804_ u2.mem\[11\]\[2\] _03857_ _03860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_165_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07529_ _02997_ _02998_ _02999_ _03000_ _03001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_74_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07598__I _02579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06277__B2 u2.mem\[155\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10540_ _05090_ _00911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10471_ _05050_ _05051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_12210_ _00089_ clknet_leaf_232_clock u2.mem\[5\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13190_ _01069_ clknet_leaf_279_clock u2.mem\[135\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07777__A1 _03229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12141_ _00020_ clknet_leaf_211_clock u2.mem\[1\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10620__I1 u2.mem\[58\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12072_ data_in_trans\[11\].A clknet_leaf_28_clock data_in_trans\[11\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11023_ _05393_ _01091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06737__C1 u2.mem\[145\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06752__A2 _02155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10136__I0 _04786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12974_ _00853_ clknet_leaf_261_clock u2.mem\[53\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12637__CLK clknet_leaf_192_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11925_ _05956_ _01430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11856_ _03679_ _05915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10807_ _05256_ _01012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09454__A1 _04417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11787_ _03670_ _05872_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08501__I0 _03811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12787__CLK clknet_leaf_26_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13526_ _01405_ clknet_leaf_314_clock u2.mem\[191\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10738_ _05195_ _05214_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_140_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12066__D data_in_trans\[8\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08009__A2 _03461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13457_ _01336_ clknet_leaf_304_clock u2.mem\[179\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10669_ _05170_ _00960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12017__CLK clknet_2_2__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12408_ _00287_ clknet_leaf_122_clock u2.mem\[17\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07217__B1 _02665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11939__I1 u2.mem\[193\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08333__S _03694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13388_ _01267_ clknet_leaf_355_clock u2.mem\[168\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07768__B2 u2.mem\[24\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12339_ _00218_ clknet_leaf_77_clock u2.mem\[13\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10611__I1 u2.mem\[58\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_290_clock_I clknet_5_20_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06440__A1 _01809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06440__B2 _01937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08568__I0 _03831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12167__CLK clknet_leaf_109_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06991__A2 _02467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06900_ _01984_ _02009_ _02379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07880_ _03342_ _03343_ _03344_ _03345_ _03346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__13412__CLK clknet_leaf_344_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06728__C1 u2.mem\[181\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06831_ u2.mem\[155\]\[5\] _02029_ _02034_ u2.mem\[174\]\[5\] u2.mem\[181\]\[5\]
+ _02038_ _02311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_23_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09550_ _04476_ u2.mem\[33\]\[5\] _04474_ _04477_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10103__S _04820_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06762_ u2.mem\[166\]\[3\] _02097_ _02099_ u2.mem\[161\]\[3\] _02243_ _02244_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08501_ _03811_ u2.mem\[9\]\[5\] _03809_ _03812_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13562__CLK clknet_leaf_40_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09481_ _04433_ _00509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06693_ _02105_ _02177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08740__I0 _03939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08432_ _03768_ _00125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08363_ _03658_ _03726_ _03633_ _03727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__10837__I mem_address_trans\[6\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07314_ _02435_ _02789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08294_ _03670_ _03671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07245_ u2.mem\[29\]\[2\] _02565_ _02570_ u2.mem\[11\]\[2\] _02722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07176_ _02520_ _02654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06127_ _01549_ _01585_ _01634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10572__I _03691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09138__I _04202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06431__A1 _01727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06058_ _01557_ _01561_ _01564_ _01565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_160_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08559__I0 _03822_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13092__CLK clknet_leaf_24_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10366__I0 _04913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09817_ _04586_ u2.mem\[39\]\[6\] _04644_ _04647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06734__A2 _02174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07931__B2 u2.mem\[62\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10013__S _04762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09748_ data_in_trans\[12\].data_sync _04604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09679_ _04482_ u2.mem\[36\]\[8\] _04554_ _04555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08731__I0 _03930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11710_ _05823_ _01348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12690_ _00569_ clknet_5_27_0_clock u2.mem\[35\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07695__B1 _03022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06498__B2 _01980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11641_ _05781_ _01321_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11618__I0 _05758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11572_ _05411_ _05729_ _05738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_167_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13311_ _01190_ clknet_leaf_347_clock u2.mem\[155\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11779__S _05866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10523_ _05007_ u2.mem\[56\]\[6\] _05078_ _05081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput19 data_in_a[6] net19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09249__S _04290_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13242_ _01121_ clknet_leaf_278_clock u2.mem\[143\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06670__A1 _02108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10454_ _05041_ _00874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08798__I0 _03917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13173_ _01052_ clknet_leaf_263_clock u2.mem\[132\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13435__CLK clknet_leaf_350_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10385_ _04994_ _04995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12124_ _01465_ clknet_leaf_36_clock u2.driver_mem\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_12_clock_I clknet_5_3_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12055_ net16 clknet_2_2__leaf_clock_a data_in_trans\[3\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10357__I0 _04904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07791__I _02456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11006_ _05381_ _05382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_42_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11019__S _05381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09712__S _04567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11857__I0 _05915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12957_ _00836_ clknet_leaf_196_clock u2.mem\[52\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10858__S _05287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08722__I0 _03921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07686__B1 _03089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_237_clock_I clknet_5_19_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11908_ _05946_ _01423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08328__S _03694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12888_ _00767_ clknet_leaf_57_clock u2.mem\[47\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11839_ _03655_ _05903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08127__I _03518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13509_ _01388_ clknet_leaf_335_clock u2.mem\[188\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07453__A3 _02919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07030_ _02508_ _02509_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_173_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06870__I _02348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08789__I0 _03908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10392__I _04138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09450__I1 u2.mem\[30\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10596__I0 _05128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08981_ _04110_ _00332_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12802__CLK clknet_leaf_145_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07932_ u2.mem\[37\]\[14\] _03291_ _03292_ u2.mem\[59\]\[14\] _03397_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10348__I0 _04895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07863_ _03320_ _03323_ _03326_ _03329_ _03330_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08705__A3 _03878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07913__A1 _03374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09602_ _04510_ _00553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06814_ u2.mem\[169\]\[4\] _02142_ _02144_ u2.mem\[147\]\[4\] _02294_ _02295_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_95_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12952__CLK clknet_leaf_49_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07794_ _02464_ _03261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09533_ _04464_ _04465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06745_ u2.mem\[153\]\[2\] _02196_ _02200_ u2.mem\[160\]\[2\] _02228_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11848__I0 _05909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11951__I _05970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08713__I0 _03912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09464_ _04418_ _04424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_149_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06676_ u2.mem\[169\]\[0\] _02142_ _02144_ u2.mem\[147\]\[0\] _02160_ _02161_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07141__A2 _02617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08415_ _03753_ _03759_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_36_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09395_ _04380_ u2.mem\[29\]\[10\] _04376_ _04381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09269__I1 u2.mem\[26\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08346_ data_in_trans\[13\].data_sync _03713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08037__I _03496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12332__CLK clknet_leaf_206_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08277_ _03656_ _03657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13458__CLK clknet_leaf_306_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07228_ u2.mem\[50\]\[2\] _02645_ _02646_ u2.mem\[51\]\[2\] _02705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06652__A1 _02006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07159_ u2.mem\[40\]\[1\] _02406_ _02415_ u2.mem\[30\]\[1\] _02637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_156_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10587__I0 _05121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09441__I1 u2.mem\[30\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06404__A1 u2.mem\[146\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12482__CLK clknet_leaf_164_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06404__B2 u2.mem\[186\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10170_ _03478_ _03986_ _04861_ _04862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_154_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06955__A2 _02391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_186_clock_I clknet_5_31_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10339__I0 _04885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08500__I _03680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07904__A1 u2.mem\[8\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06707__A2 _02030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08952__I0 _04048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07904__B2 u2.mem\[4\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12811_ _00690_ clknet_leaf_221_clock u2.mem\[43\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12742_ _00621_ clknet_leaf_70_clock u2.mem\[38\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12673_ _00552_ clknet_leaf_154_clock u2.mem\[34\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11624_ _05746_ u2.mem\[176\]\[0\] _05771_ _05772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11555_ _05719_ u2.mem\[171\]\[5\] _05721_ _05728_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06643__A1 _02108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10506_ _05070_ _00897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11486_ _05671_ u2.mem\[167\]\[2\] _05683_ _05686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12825__CLK clknet_leaf_136_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13225_ _01104_ clknet_leaf_283_clock u2.mem\[141\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10437_ _04992_ u2.mem\[54\]\[1\] _05030_ _05032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07199__A2 _02580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13156_ _01035_ clknet_leaf_262_clock u2.mem\[129\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10368_ _04916_ u2.mem\[52\]\[13\] _04981_ _04983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12107_ _01490_ clknet_leaf_135_clock u2.active_mem\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10940__I _04126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13087_ _00966_ clknet_leaf_245_clock u2.mem\[60\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12975__CLK clknet_leaf_249_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10299_ _04072_ _04863_ _04943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09196__I0 _04254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12038_ col_select_trans\[0\].A clknet_leaf_302_clock col_select_trans\[0\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08943__I0 _04039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12205__CLK clknet_leaf_212_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07026__I _02504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06530_ _01998_ _02015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07659__B1 _03050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06461_ u2.mem\[0\]\[8\] _01954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12355__CLK clknet_leaf_83_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08200_ _03548_ u2.mem\[3\]\[1\] _03609_ _03611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09180_ _04171_ u2.mem\[24\]\[13\] _04241_ _04243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06392_ _01891_ _01892_ _01893_ _01894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_1565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08131_ _03521_ _03566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08062_ _03515_ _03508_ _03516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07831__B1 _03140_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07013_ _02432_ _02492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_128_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06105__I _01561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08964_ _04021_ u2.mem\[20\]\[3\] _04097_ _04101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09416__I _04395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07915_ u2.mem\[1\]\[14\] _03261_ _03262_ u2.mem\[7\]\[14\] _03380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08320__I _03691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08895_ _04030_ u2.mem\[18\]\[7\] _04056_ _04060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08934__I0 _04030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_341_clock clknet_5_5_0_clock clknet_leaf_341_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_5_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07846_ _02600_ _03313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_5_20_0_clock_I clknet_4_10_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06165__A3 _01582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input17_I data_in_a[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13130__CLK clknet_leaf_327_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07777_ _03229_ _03234_ _03239_ _03244_ _03245_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_99_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09516_ _04378_ u2.mem\[32\]\[9\] _04453_ _04455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06728_ u2.mem\[155\]\[2\] _02030_ _02035_ u2.mem\[174\]\[2\] u2.mem\[181\]\[2\]
+ _02039_ _02211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_38_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_356_clock clknet_5_1_0_clock clknet_leaf_356_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_38_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08162__I1 u2.mem\[2\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09447_ _04413_ _00495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_06659_ _02143_ _02144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13280__CLK clknet_leaf_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09378_ _04144_ _04369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12848__CLK clknet_leaf_151_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08329_ _03699_ _00091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11122__S _05453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11340_ _05592_ _01209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06625__A1 u2.mem\[159\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06625__B2 u2.mem\[149\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06443__C _01934_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11271_ _05549_ _01183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13010_ _00889_ clknet_leaf_237_clock u2.mem\[55\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_165_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09527__S _04458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10222_ _04894_ _00789_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06389__B1 _01635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11856__I _03679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10153_ _04852_ _00762_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09178__I0 _04167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12228__CLK clknet_leaf_64_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10980__I0 _05340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10084_ _04810_ u2.mem\[45\]\[12\] _04811_ _04812_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09878__A1 _04249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_309_clock clknet_5_16_0_clock clknet_leaf_309_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08925__I0 _04021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11685__A1 _04094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10732__I0 _05209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09262__S _04295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12378__CLK clknet_leaf_60_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11591__I _05667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10201__S _04880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11288__I1 u2.mem\[155\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10986_ _05349_ u2.mem\[136\]\[4\] _05364_ _05370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12725_ _00604_ clknet_leaf_72_clock u2.mem\[37\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12656_ _00535_ clknet_leaf_221_clock u2.mem\[33\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09102__I0 _04167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10935__I _05334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11607_ _05760_ _05761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_12587_ _00466_ clknet_leaf_186_clock u2.mem\[29\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09802__A1 _03752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11032__S _05395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06616__A1 _01992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07813__B1 _03124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11538_ _05717_ u2.mem\[170\]\[4\] _05708_ _05718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11967__S _05980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12074__D data_in_trans\[12\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13003__CLK clknet_leaf_249_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11469_ _05673_ _05674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09437__S _04406_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13208_ _01087_ clknet_leaf_281_clock u2.mem\[138\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07041__A1 _02394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13139_ _01018_ clknet_leaf_21_clock u2.mem\[63\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10971__I0 _05349_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09169__I0 _04154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input9_I data_in_a[11] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13153__CLK clknet_leaf_268_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08140__I _03528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07700_ u2.mem\[3\]\[10\] _03034_ _02978_ _03169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_152_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08680_ _03905_ _03924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_22_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07631_ u2.mem\[45\]\[9\] _03099_ _03100_ u2.mem\[34\]\[9\] _03101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11207__S _05502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07562_ u2.mem\[16\]\[8\] _03031_ _03032_ u2.mem\[33\]\[8\] _03033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11279__I1 u2.mem\[154\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09301_ _04267_ u2.mem\[27\]\[7\] _04318_ _04322_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06513_ row_select_trans\[5\].data_sync _01997_ _01998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07493_ u2.mem\[8\]\[6\] _02858_ _02859_ u2.mem\[4\]\[6\] _02966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_134_clock_I clknet_5_12_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11006__I _05381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09232_ _04278_ u2.mem\[25\]\[12\] _04279_ _04280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06444_ _01844_ _01938_ _01939_ _01940_ _01468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_61_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06855__B2 u2.mem\[147\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09163_ _04233_ _00391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06375_ u2.mem\[0\]\[5\] _01877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_33_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08114_ _03507_ _03554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09094_ _04193_ _00362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08315__I _03687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07804__B1 _03115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08045_ _03502_ _03503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07280__B2 u2.mem\[20\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09347__S _04346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11203__I1 u2.mem\[150\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09996_ _04709_ u2.mem\[43\]\[12\] _04755_ _04756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_280_clock clknet_5_21_0_clock clknet_leaf_280_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07583__A2 _02899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_59_clock_I clknet_5_12_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08050__I _03506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08947_ _04090_ _00318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06791__B1 _02244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08907__I0 _04041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12520__CLK clknet_leaf_118_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08878_ _03583_ _03988_ _04050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_3826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06138__A3 _01600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07829_ u2.mem\[57\]\[12\] _03294_ _03295_ u2.mem\[41\]\[12\] _03296_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_3859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07886__A3 _03346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_295_clock clknet_5_17_0_clock clknet_leaf_295_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_56_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10840_ _05275_ _05276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_77_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09810__S _04639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10771_ _05202_ u2.mem\[62\]\[3\] _05232_ _05236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12510_ _00389_ clknet_leaf_179_clock u2.mem\[24\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06846__A1 u2.mem\[153\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13490_ _01369_ clknet_leaf_292_clock u2.mem\[185\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12441_ _00320_ clknet_leaf_127_clock u2.mem\[19\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13026__CLK clknet_leaf_251_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12372_ _00251_ clknet_leaf_80_clock u2.mem\[15\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11442__I1 u2.mem\[165\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_233_clock clknet_5_18_0_clock clknet_leaf_233_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_165_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11323_ _05554_ u2.mem\[157\]\[4\] _05575_ _05581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_336_clock_I clknet_5_4_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11254_ _05505_ u2.mem\[153\]\[1\] _05537_ _05539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10205_ _04815_ u2.mem\[48\]\[14\] _04880_ _04883_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07023__A1 _02483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11185_ _05464_ u2.mem\[149\]\[1\] _05492_ _05494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_248_clock clknet_5_22_0_clock clknet_leaf_248_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09056__I _04123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07574__A2 _03038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10136_ _04786_ u2.mem\[47\]\[1\] _04841_ _04843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06782__B1 _02019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10067_ _04799_ u2.mem\[45\]\[7\] _04793_ _04800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12069__D net8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10866__S _05286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08826__A2 _04013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11130__I0 _05432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10969_ _05346_ u2.mem\[135\]\[3\] _05356_ _05360_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06837__A1 u2.mem\[159\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12708_ _00587_ clknet_leaf_68_clock u2.mem\[36\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06837__B2 u2.mem\[149\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12639_ _00518_ clknet_leaf_175_clock u2.mem\[32\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06160_ _01666_ _01667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13519__CLK clknet_leaf_16_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11697__S _05809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06065__A2 _01571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07262__B2 u2.mem\[2\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06091_ u2.mem\[166\]\[0\] _01592_ _01595_ u2.mem\[149\]\[0\] _01597_ u2.mem\[161\]\[0\]
+ _01598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_144_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11496__I _05691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12543__CLK clknet_leaf_168_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07014__A1 _02401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09850_ _04660_ _04666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10106__S _04825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08801_ _03998_ _00264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_60_clock_I clknet_5_12_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_06993_ u2.mem\[1\]\[0\] _02465_ _02471_ u2.mem\[7\]\[0\] _02472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09781_ _04626_ _00616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08732_ _03956_ _00237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08663_ _03671_ _03912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07614_ u2.mem\[18\]\[8\] _03083_ _03084_ u2.mem\[19\]\[8\] _03085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08594_ _03820_ u2.mem\[11\]\[9\] _03867_ _03869_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07545_ _02395_ _03016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10776__S _05237_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_12_0_clock clknet_3_6_0_clock clknet_4_12_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_clkbuf_leaf_285_clock_I clknet_5_20_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06828__A1 u2.mem\[184\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07476_ u2.mem\[61\]\[6\] _02899_ _02900_ u2.mem\[63\]\[6\] _02949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08246__S _03635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11672__I1 u2.mem\[179\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09215_ _04267_ u2.mem\[25\]\[7\] _04261_ _04268_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06427_ _01916_ _01927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06274__B _01554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09146_ _04222_ _00385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12073__CLK clknet_2_1__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13199__CLK clknet_leaf_274_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06358_ u2.mem\[166\]\[4\] _01753_ _01754_ u2.mem\[161\]\[4\] _01860_ _01861_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08045__I _03502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06056__A2 col_select_trans\[1\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09077_ _04128_ u2.mem\[22\]\[1\] _04182_ _04184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06289_ u2.mem\[190\]\[2\] _01703_ _01705_ u2.mem\[194\]\[2\] _01794_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11400__S _05625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09077__S _04182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08028_ _03488_ _03489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07005__A1 _02440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10016__S _04767_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09979_ _04746_ _00694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07020__A4 _02498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12990_ _00869_ clknet_leaf_258_clock u2.mem\[54\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09553__I0 _04478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11941_ _05949_ _05965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_3645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11872_ _05924_ _01409_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07124__I _02602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09540__S _04465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10686__S _05179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10823_ _05265_ _01019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11112__I0 _05428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06819__A1 u2.mem\[154\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06819__B2 u2.mem\[162\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13542_ _01421_ clknet_leaf_21_clock u2.mem\[192\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10754_ _03713_ _05225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13473_ _01352_ clknet_leaf_292_clock u2.mem\[182\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10685_ _05180_ _00966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_172_clock clknet_5_27_0_clock clknet_leaf_172_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_145_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12424_ _00303_ clknet_leaf_123_clock u2.mem\[18\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11415__I1 u2.mem\[163\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07244__A1 u2.mem\[26\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12566__CLK clknet_leaf_94_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12355_ _00234_ clknet_leaf_83_clock u2.mem\[14\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07794__I _02464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11306_ _05571_ _01196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12286_ _00165_ clknet_leaf_185_clock u2.mem\[10\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11179__I0 _05472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_187_clock clknet_5_31_0_clock clknet_leaf_187_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_153_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11237_ _05528_ _05529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_106_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10926__I0 _05301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06203__I _01709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11168_ _05483_ _05484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_68_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_110_clock clknet_5_14_0_clock clknet_leaf_110_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10119_ _04806_ u2.mem\[46\]\[10\] _04830_ _04833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11099_ _05440_ _01120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11351__I0 _05587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11980__S _05985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_125_clock clknet_5_15_0_clock clknet_leaf_125_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_17_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07330_ u2.mem\[54\]\[4\] _02648_ _02649_ u2.mem\[55\]\[4\] _02805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12096__CLK clknet_leaf_214_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13341__CLK clknet_leaf_3_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07483__A1 u2.mem\[9\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07261_ u2.mem\[45\]\[3\] _02633_ _02634_ u2.mem\[34\]\[3\] _02737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06286__A2 _01565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09000_ _04123_ _04124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12909__CLK clknet_leaf_202_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06212_ _01612_ _01613_ _01596_ _01719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_136_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06691__C1 u2.mem\[159\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11406__I1 u2.mem\[162\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07192_ u2.mem\[37\]\[1\] _02540_ _02542_ u2.mem\[59\]\[1\] _02670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_157_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06143_ _01649_ _01650_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13491__CLK clknet_leaf_292_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10090__I0 _04815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06074_ _01580_ _01581_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09902_ _04698_ u2.mem\[41\]\[7\] _04692_ _04699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07209__I _02626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09625__S _04522_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09833_ _04609_ u2.mem\[39\]\[13\] _04654_ _04656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06746__B1 _02130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09764_ _04616_ _00609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_06976_ _02454_ _02455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_100_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08715_ _03941_ _03947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_55_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10145__I1 u2.mem\[47\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09695_ _04563_ _00593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11342__I0 _05593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08646_ _03833_ u2.mem\[12\]\[15\] _03895_ _03899_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_76_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12439__CLK clknet_leaf_127_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07710__A2 _03049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08577_ _03859_ _00179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07528_ u2.mem\[28\]\[7\] _02839_ _02840_ u2.mem\[31\]\[7\] _03000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07069__A4 _02411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07459_ _02928_ _02929_ _02930_ _02931_ _02932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_126_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12589__CLK clknet_leaf_187_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10470_ _03752_ _04964_ _05050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06029__A2 _01517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09129_ _04202_ _04213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_100_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07777__A2 _03234_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12140_ _00019_ clknet_leaf_211_clock u2.mem\[1\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08503__I _03684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12071_ net9 clknet_2_1__leaf_clock_a data_in_trans\[11\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10908__I0 _05294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07119__I _02597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11022_ _05392_ u2.mem\[138\]\[5\] _05381_ _05393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06737__C2 _02081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12973_ _00852_ clknet_leaf_262_clock u2.mem\[53\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11333__I0 _05587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_42_clock clknet_5_6_0_clock clknet_leaf_42_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_4187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11924_ _05913_ u2.mem\[193\]\[4\] _05955_ _05956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07162__B1 _02461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13364__CLK clknet_leaf_358_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11855_ _05914_ _01402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11305__S _05568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06693__I _02105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10806_ u2.mem\[63\]\[2\] _03500_ _05253_ _05256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_57_clock clknet_5_12_0_clock clknet_leaf_57_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_14_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11786_ _05871_ _01376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08501__I1 u2.mem\[9\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13525_ _01404_ clknet_leaf_315_clock u2.mem\[191\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10737_ _03691_ _05213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13456_ _01335_ clknet_leaf_304_clock u2.mem\[179\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10668_ _05126_ u2.mem\[59\]\[14\] _05167_ _05170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12407_ _00286_ clknet_leaf_112_clock u2.mem\[17\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07217__A1 _01726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13387_ _01266_ clknet_leaf_355_clock u2.mem\[168\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10599_ _05130_ _05131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_127_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07768__A2 _03077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12338_ _00217_ clknet_leaf_152_clock u2.mem\[13\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_233_clock_I clknet_5_18_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06440__A2 _01915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12269_ _00148_ clknet_leaf_185_clock u2.mem\[9\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08568__I1 u2.mem\[10\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06830_ u2.mem\[150\]\[5\] _02192_ _02310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06868__I _02346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09244__I _04287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07940__A2 _02596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06761_ _02240_ _02241_ _02242_ _02243_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_55_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08500_ _03680_ _03811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09480_ _04382_ u2.mem\[31\]\[11\] _04429_ _04433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06692_ _02109_ _02176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08740__I1 u2.mem\[14\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08431_ _03706_ u2.mem\[7\]\[11\] _03764_ _03768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12731__CLK clknet_leaf_216_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11215__S _05501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08362_ _03725_ _03606_ _03726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_36_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07313_ _02427_ _02788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07456__A1 u2.mem\[32\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08293_ _03502_ _03670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07244_ u2.mem\[26\]\[2\] _02673_ _02674_ u2.mem\[10\]\[2\] _02721_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12881__CLK clknet_leaf_143_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07175_ _02647_ _02650_ _02651_ _02652_ _02653_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_118_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08956__A1 _04095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06126_ _01632_ _01633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10763__A1 _04394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11885__S _05932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12111__CLK clknet_leaf_332_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06057_ _01563_ _01564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06431__A2 _01915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10366__I1 u2.mem\[52\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11684__I _05768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09816_ _04646_ _00631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06195__A1 _01561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12261__CLK clknet_leaf_70_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13387__CLK clknet_leaf_355_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09747_ _04603_ _00605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06959_ _02370_ _02438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__11315__I0 _05544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09678_ _04543_ _04554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_36_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08731__I1 u2.mem\[14\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07695__A1 u2.mem\[27\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08629_ _03889_ _00201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06498__A2 _01924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11640_ _05750_ u2.mem\[177\]\[1\] _05779_ _05781_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_182_clock_I clknet_5_27_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11571_ _05737_ _01295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13310_ _01189_ clknet_leaf_348_clock u2.mem\[155\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10522_ _05080_ _00903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08434__S _03769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13241_ _01120_ clknet_leaf_272_clock u2.mem\[143\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10453_ _05011_ u2.mem\[54\]\[8\] _05040_ _05041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06670__A2 _02052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10054__I0 _04790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13172_ _01051_ clknet_leaf_263_clock u2.mem\[132\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10384_ _04130_ _04994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06958__B1 _02436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12123_ _01458_ clknet_leaf_37_clock u2.driver_mem\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09265__S _04300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12054_ data_in_trans\[2\].A clknet_leaf_287_clock data_in_trans\[2\].data_sync vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11005_ _04288_ _05363_ _05381_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_46_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06186__A1 _01563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09064__I _04173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12956_ _00835_ clknet_leaf_197_clock u2.mem\[52\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_1574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11857__I1 u2.mem\[190\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08722__I1 u2.mem\[14\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11907_ u2.mem\[192\]\[13\] _03531_ _05942_ _05946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12887_ _00766_ clknet_leaf_57_clock u2.mem\[47\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11838_ _05902_ _01397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12077__D net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10874__S _05297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11769_ _05860_ _01370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10293__I0 _04916_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13508_ _01387_ clknet_leaf_331_clock u2.mem\[188\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08344__S _03711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07453__A4 _02926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12134__CLK clknet_leaf_14_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13439_ _01318_ clknet_leaf_341_clock u2.mem\[176\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10045__I0 _04782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08980_ _04037_ u2.mem\[20\]\[10\] _04107_ _04110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12284__CLK clknet_leaf_185_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09175__S _04236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09738__I0 _04596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07931_ u2.mem\[60\]\[14\] _03288_ _03289_ u2.mem\[62\]\[14\] _03396_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_155_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11545__I0 _05707_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07862_ u2.mem\[6\]\[12\] _03327_ _03328_ u2.mem\[47\]\[12\] _03329_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09601_ _04480_ u2.mem\[34\]\[7\] _04506_ _04510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06813_ _02291_ _02292_ _02293_ _02294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07793_ u2.mem\[15\]\[12\] _03258_ _03259_ u2.mem\[13\]\[12\] _03260_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11009__I _05339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09532_ _04013_ _04441_ _04464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_83_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06744_ u2.mem\[194\]\[2\] _02198_ _02199_ u2.mem\[190\]\[2\] _02227_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11848__I1 u2.mem\[190\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09702__I _04126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09463_ _04423_ _00501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06675_ _02149_ _02154_ _02159_ _02160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08414_ _03758_ _00117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09394_ _04160_ _04380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08345_ _03712_ _00094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10284__I0 _04907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08276_ _03655_ _03656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08229__I0 _03577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07227_ _02700_ _02701_ _02702_ _02703_ _02704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06652__A2 _02002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10036__I0 _04712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07158_ u2.mem\[32\]\[1\] _02386_ _02396_ u2.mem\[2\]\[1\] _02636_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12627__CLK clknet_leaf_97_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06109_ _01580_ _01616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06404__A2 _01691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07089_ _02363_ _02568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_65_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09729__I0 _04589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06955__A3 _02424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_129_clock_I clknet_5_14_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10339__I1 u2.mem\[52\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12777__CLK clknet_leaf_130_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06168__A1 _01638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12810_ _00689_ clknet_leaf_139_clock u2.mem\[42\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12007__CLK clknet_2_2__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09612__I _04500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12741_ _00620_ clknet_leaf_70_clock u2.mem\[38\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07668__A1 _03134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12672_ _00551_ clknet_leaf_177_clock u2.mem\[34\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12157__CLK clknet_leaf_205_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11623_ _05770_ _05771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13402__CLK clknet_leaf_298_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10275__I0 _04898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08093__A1 u2.driver_enable vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08164__S _03585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11554_ _05727_ _01288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_1458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10505_ _05027_ u2.mem\[55\]\[15\] _05066_ _05070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06643__A2 _02041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11485_ _05685_ _01261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10027__I0 _04703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09059__I data_in_trans\[13\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13224_ _01103_ clknet_leaf_286_clock u2.mem\[140\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10436_ _05031_ _00866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08640__I0 _03826_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13155_ _01034_ clknet_leaf_261_clock u2.mem\[129\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10367_ _04982_ _00846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12106_ _01489_ clknet_leaf_58_clock u2.active_mem\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06946__A3 _02424_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13086_ _00965_ clknet_leaf_267_clock u2.mem\[60\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10298_ _04942_ _00817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12037_ net1 clknet_2_0__leaf_clock_a col_select_trans\[0\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06159__A1 _01638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11152__A1 _04071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07307__I _02385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08943__I1 u2.mem\[19\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09522__I _04442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07659__B2 u2.mem\[20\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12939_ _00818_ clknet_leaf_251_clock u2.mem\[51\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06460_ _01951_ _01938_ _01952_ _01953_ _01471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_61_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06331__A1 u2.mem\[173\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07042__I _02520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06331__B2 u2.mem\[185\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06391_ u2.mem\[159\]\[5\] _01603_ _01594_ u2.mem\[149\]\[5\] _01893_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13082__CLK clknet_leaf_42_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08130_ _03565_ _00026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10266__I0 _04889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06881__I _02359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08084__A1 _03531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08061_ data_in_trans\[7\].data_sync _03515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_174_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07831__B2 u2.mem\[10\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10018__I0 _04694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07012_ _02430_ _02491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_134_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09959__I0 _04709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08802__S _03995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11766__I0 _05829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09584__A1 _03583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08631__I0 _03817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_130_clock_I clknet_5_14_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08963_ _04100_ _00324_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07914_ u2.mem\[15\]\[14\] _03258_ _03259_ u2.mem\[13\]\[14\] _03379_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08894_ _04059_ _00296_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08934__I1 u2.mem\[19\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07845_ u2.mem\[17\]\[12\] _03310_ _03311_ u2.mem\[24\]\[12\] _03312_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07776_ _03240_ _03241_ _03242_ _03243_ _03244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_77_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09515_ _04454_ _00522_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06727_ u2.mem\[150\]\[2\] _02192_ _02210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_24_0_clock_I clknet_4_12_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13425__CLK clknet_leaf_349_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09446_ _04387_ u2.mem\[30\]\[13\] _04411_ _04413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08048__I _03489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06658_ _02023_ _02077_ _02143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09377_ _04368_ _00470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06589_ _02056_ _02063_ _02069_ _02073_ _02074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_138_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_55_clock_I clknet_5_12_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11403__S _05625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10257__I0 _04918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08328_ _03698_ u2.mem\[5\]\[9\] _03694_ _03699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13575__CLK clknet_leaf_34_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08870__I0 _04044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08259_ _03646_ _00074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10009__I0 _04685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11202__I _05504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09808__S _04639_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11270_ _05548_ u2.mem\[154\]\[1\] _05546_ _05549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10221_ _04893_ u2.mem\[49\]\[3\] _04887_ _04894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08622__I0 _03808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06389__A1 u2.mem\[187\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06389__B2 u2.mem\[192\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07586__B1 _03056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10152_ _04801_ u2.mem\[47\]\[8\] _04851_ _04852_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07050__A2 _02526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10083_ _04783_ _04811_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07338__B1 _02655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07127__I _02605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09543__S _04465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09878__A2 _04659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11685__A2 _05808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10732__I1 u2.mem\[61\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06966__I _02430_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09342__I _04335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_332_clock_I clknet_5_7_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10985_ _05369_ _01077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10496__I0 _05018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12724_ _00603_ clknet_leaf_72_clock u2.mem\[37\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06313__A1 u2.mem\[189\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07510__B1 _02882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12655_ _00534_ clknet_leaf_223_clock u2.mem\[33\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07797__I _02474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09102__I1 u2.mem\[22\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11606_ _04416_ _05729_ _05760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_12586_ _00465_ clknet_leaf_115_clock u2.mem\[28\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07813__A1 u2.mem\[14\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11537_ _05676_ _05717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06616__A2 _02002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07813__B2 u2.mem\[12\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06206__I _01712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08622__S _03885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11468_ _03502_ _05673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13207_ _01086_ clknet_leaf_287_clock u2.mem\[138\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08613__I0 _03798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10419_ _05019_ _00861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07577__B1 _02894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11399_ _05507_ _05629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13138_ _01017_ clknet_leaf_314_clock u2.mem\[63\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13069_ _00948_ clknet_leaf_259_clock u2.mem\[59\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07329__B1 _02646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12322__CLK clknet_leaf_158_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13448__CLK clknet_leaf_343_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07630_ _02447_ _03100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07561_ _02476_ _03032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10398__I _05004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09300_ _04321_ _00440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06512_ row_select_trans\[4\].data_sync _01997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10487__I0 _05009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07492_ u2.mem\[39\]\[6\] _02855_ _02856_ u2.mem\[48\]\[6\] _02965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12472__CLK clknet_leaf_121_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09231_ _04251_ _04279_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_146_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06855__A2 _02141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06443_ u2.mem\[193\]\[4\] _01928_ _01929_ u2.mem\[192\]\[4\] _01934_ _01940_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_167_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11223__S _05520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09162_ _04145_ u2.mem\[24\]\[5\] _04231_ _04233_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06374_ _01844_ _01555_ _01876_ _01484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08057__A1 _01878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08113_ _03553_ _00021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09093_ _04154_ u2.mem\[22\]\[8\] _04192_ _04193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08044_ data_in_trans\[3\].data_sync _03502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07280__A2 _02515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11739__I0 _05831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11957__I _05971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08331__I _03700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_281_clock_I clknet_5_21_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09995_ _04739_ _04755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_88_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08946_ _04041_ u2.mem\[19\]\[12\] _04089_ _04090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06791__A1 _01809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09363__S _04358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06791__B2 _02272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08877_ _04049_ _00289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07828_ _02555_ _03295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07886__A4 _03351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07759_ u2.mem\[37\]\[11\] _03058_ _03059_ u2.mem\[59\]\[11\] _03227_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10478__I0 _04998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10770_ _05235_ _00996_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08707__S _03942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09429_ _04403_ _00487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06846__A2 _02136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12965__CLK clknet_leaf_85_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12440_ _00319_ clknet_leaf_123_clock u2.mem\[19\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08506__I _03688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11978__I0 _05220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12371_ _00250_ clknet_leaf_78_clock u2.mem\[15\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11322_ _05580_ _01203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10650__I0 _05108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07271__A2 _02743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11253_ _05538_ _01176_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07559__B1 _03029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10204_ _04882_ _00783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10402__I0 _05007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11184_ _05493_ _01152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12345__CLK clknet_leaf_60_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10135_ _04842_ _00754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06782__B2 u2.mem\[189\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10066_ _04588_ _04799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10212__S _04887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06534__A1 _02015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12495__CLK clknet_leaf_163_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07731__B1 _03095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09072__I _04179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08617__S _03880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10968_ _05359_ _01070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11130__I1 u2.mem\[145\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12707_ _00586_ clknet_leaf_30_clock u2.mem\[36\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11043__S _05404_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10899_ _05303_ u2.mem\[131\]\[3\] _05310_ _05314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08039__A1 _01727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12638_ _00517_ clknet_leaf_192_clock u2.mem\[32\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07320__I _02464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06364__C _01866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11969__I0 _05211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12085__D net34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11978__S _05985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_340_clock clknet_5_5_0_clock clknet_leaf_340_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12569_ _00448_ clknet_leaf_113_clock u2.mem\[27\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08834__I0 _04019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10641__I0 _05099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06090_ _01576_ _01596_ _01597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_172_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_355_clock clknet_5_1_0_clock clknet_leaf_355_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07014__A2 _02403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08800_ _03919_ u2.mem\[16\]\[6\] _03995_ _03998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13270__CLK clknet_leaf_5_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09780_ _04586_ u2.mem\[38\]\[6\] _04623_ _04626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06992_ _02470_ _02471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08731_ _03930_ u2.mem\[14\]\[11\] _03952_ _03956_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12838__CLK clknet_leaf_63_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09011__I0 _04132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08662_ _03911_ _00212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07613_ _02607_ _03084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08593_ _03868_ _00186_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12988__CLK clknet_leaf_257_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07544_ _02385_ _03015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_228_clock_I clknet_5_25_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09710__I _04134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06289__B1 _01705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07475_ _02932_ _02937_ _02942_ _02947_ _02948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_22_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09214_ _04150_ _04267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12218__CLK clknet_leaf_52_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10880__I0 _05301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06426_ u2.mem\[194\]\[1\] _01924_ _01926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08326__I _03696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09145_ _04177_ u2.mem\[23\]\[15\] _04218_ _04222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06357_ _01857_ _01858_ _01859_ _01860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_108_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09076_ _04183_ _00354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08262__S _03645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06288_ _01789_ _01790_ _01791_ _01792_ _01793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_11_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08027_ _03480_ _03487_ _03488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07005__A2 _02441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08061__I data_in_trans\[7\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09978_ _04691_ u2.mem\[43\]\[4\] _04745_ _04746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06764__A1 u2.mem\[194\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09093__S _04192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06764__B2 u2.mem\[190\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08929_ _04080_ _00310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10699__I0 _05119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09553__I1 u2.mem\[33\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11940_ _05964_ _01437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07405__I _02504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07713__B1 _03133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10967__S _05356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11871_ _05915_ u2.mem\[191\]\[5\] _05917_ _05924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10822_ u2.mem\[63\]\[9\] _03521_ _05263_ _05265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11112__I1 u2.mem\[144\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13541_ _01420_ clknet_leaf_21_clock u2.mem\[192\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10753_ _05224_ _00990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09069__I0 _04177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13472_ _01351_ clknet_leaf_294_clock u2.mem\[182\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10684_ _05103_ u2.mem\[60\]\[4\] _05179_ _05180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13143__CLK clknet_leaf_39_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07140__I _02618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11798__S _05879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12423_ _00302_ clknet_leaf_128_clock u2.mem\[18\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08816__I0 _03935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07244__A2 _02673_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12354_ _00233_ clknet_leaf_150_clock u2.mem\[14\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11305_ _05550_ u2.mem\[156\]\[2\] _05568_ _05571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13293__CLK clknet_leaf_364_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12285_ _00164_ clknet_leaf_185_clock u2.mem\[10\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10207__S _04880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11328__A1 _04393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09067__I data_in_trans\[15\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11236_ _04223_ _05527_ _05528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09241__I0 _04285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08900__S _04061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10006__I _04761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11167_ _04094_ _05482_ _05483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_136_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_177_clock_I clknet_5_27_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06755__A1 _02224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07952__B1 _02448_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10118_ _04832_ _00747_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11098_ _05430_ u2.mem\[143\]\[4\] _05434_ _05440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10049_ _04787_ _00723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06507__A1 row_select_trans\[5\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07704__B1 _03040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11351__I1 u2.mem\[159\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10877__S _05297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07260_ _01768_ _02361_ _02715_ _02736_ _01494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10862__I0 _05200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06140__C1 u2.mem\[165\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06211_ u2.mem\[154\]\[0\] _01699_ _01701_ u2.mem\[162\]\[0\] _01717_ _01718_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__06691__B1 _02098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07191_ u2.mem\[60\]\[1\] _02546_ _02549_ u2.mem\[62\]\[1\] _02669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08807__I0 _03926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06691__C2 _02174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12510__CLK clknet_leaf_179_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11501__S _05692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06142_ _01612_ _01616_ _01644_ _01649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__09480__I0 _04382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07235__A2 _02660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06443__B1 _01929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_294_clock clknet_5_20_0_clock clknet_leaf_294_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06073_ _01550_ _01579_ _01580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__10117__S _04830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11300__I _05567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09901_ _04588_ _04698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_160_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09232__I0 _04278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12660__CLK clknet_leaf_75_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09832_ _04655_ _00638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06746__A1 u2.mem\[148\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06746__B2 u2.mem\[152\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09763_ _04615_ u2.mem\[37\]\[15\] _04606_ _04616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06975_ _02362_ _02454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13016__CLK clknet_leaf_319_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08714_ _03946_ _00229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09694_ _04498_ u2.mem\[36\]\[15\] _04559_ _04563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09641__S _04532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11342__I1 u2.mem\[158\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08645_ _03898_ _00208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_232_clock clknet_5_24_0_clock clknet_leaf_232_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_26_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10787__S _05242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08576_ _03802_ u2.mem\[11\]\[1\] _03857_ _03859_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09299__I0 _04265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12040__CLK clknet_leaf_299_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13166__CLK clknet_leaf_263_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_07527_ u2.mem\[9\]\[7\] _02836_ _02837_ u2.mem\[25\]\[7\] _02999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_126_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10586__I _05094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10853__I0 _05207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07458_ u2.mem\[27\]\[6\] _02788_ _02789_ u2.mem\[35\]\[6\] _02931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12190__CLK clknet_leaf_252_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06409_ _01878_ _01554_ _01910_ _01485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07389_ _02854_ _02857_ _02860_ _02863_ _02864_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__11558__A1 _04333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08018__A4 mem_address_trans\[7\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09128_ _04212_ _00377_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07226__A2 _02480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09471__I0 _04373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10027__S _04772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07777__A3 _03239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09059_ data_in_trans\[13\].data_sync _04170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11210__I _05510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12070_ data_in_trans\[10\].A clknet_leaf_28_clock data_in_trans\[10\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08720__S _03947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11030__I0 _05386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11021_ _05351_ _05392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06737__A1 u2.mem\[165\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06737__B2 u2.mem\[163\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12972_ _00851_ clknet_leaf_262_clock u2.mem\[53\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07135__I _02613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11333__I1 u2.mem\[158\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11923_ _05949_ _05955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_57_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10697__S _05184_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11854_ _05913_ u2.mem\[190\]\[4\] _05904_ _05914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10805_ _05255_ _01011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11785_ _05870_ u2.mem\[186\]\[2\] _05866_ _05871_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12533__CLK clknet_leaf_98_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13524_ _01403_ clknet_leaf_15_clock u2.mem\[190\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10736_ _05212_ _00985_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13455_ _01334_ clknet_leaf_302_clock u2.mem\[179\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10667_ _05169_ _00959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11321__S _05576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12406_ _00285_ clknet_leaf_88_clock u2.mem\[17\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07217__A2 _02361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09462__I0 _04364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12683__CLK clknet_leaf_195_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13386_ _01265_ clknet_leaf_306_clock u2.mem\[167\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10598_ _04288_ _05071_ _05130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_115_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12337_ _00216_ clknet_leaf_152_clock u2.mem\[13\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12268_ _00147_ clknet_leaf_185_clock u2.mem\[9\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11219_ _05517_ u2.mem\[150\]\[5\] _05501_ _05518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12199_ _00078_ clknet_leaf_66_clock u2.mem\[4\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06728__A1 u2.mem\[155\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07925__B1 _02528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06760_ u2.mem\[188\]\[3\] _02185_ _02177_ u2.mem\[175\]\[3\] _02242_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12063__CLK clknet_2_3__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06691_ u2.mem\[166\]\[1\] _02096_ _02098_ u2.mem\[161\]\[1\] u2.mem\[159\]\[1\]
+ _02174_ _02175_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__07153__A1 _02563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11790__I _03674_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08430_ _03767_ _00124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06884__I _02362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08361_ _03481_ _03725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07312_ u2.mem\[40\]\[4\] _02785_ _02786_ u2.mem\[30\]\[4\] _02787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10835__I0 u2.mem\[63\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08653__A1 _03480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08292_ _03669_ _00084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06259__A3 _01763_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08805__S _04000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07243_ _02716_ _02717_ _02718_ _02719_ _02720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11231__S _05519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08405__A1 _03480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07174_ u2.mem\[58\]\[1\] _02495_ _02500_ u2.mem\[36\]\[1\] _02652_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11260__I0 _05514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06125_ _01616_ _01609_ _01632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09636__S _04527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06124__I _01630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06056_ _01562_ col_select_trans\[1\].data_sync _01563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_154_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09815_ _04583_ u2.mem\[39\]\[5\] _04644_ _04646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06195__A2 _01563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09746_ _04602_ u2.mem\[37\]\[11\] _04593_ _04603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_171_clock clknet_5_27_0_clock clknet_leaf_171_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06958_ u2.mem\[27\]\[0\] _02428_ _02436_ u2.mem\[35\]\[0\] _02437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11315__I1 u2.mem\[157\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09677_ _04553_ _00585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_06889_ _02353_ _02368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12556__CLK clknet_leaf_190_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11406__S _05624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08628_ _03815_ u2.mem\[12\]\[7\] _03885_ _03889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10310__S _04949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07695__A2 _03021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06352__C1 _01732_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08559_ _03822_ u2.mem\[10\]\[10\] _03846_ _03849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_186_clock clknet_5_31_0_clock clknet_leaf_186_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_125_clock_I clknet_5_15_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11205__I _03499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11570_ _05719_ u2.mem\[172\]\[5\] _05730_ _05737_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09692__I0 _04496_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06655__B1 _02127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10521_ _05005_ u2.mem\[56\]\[5\] _05078_ _05080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11141__S _05462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13240_ _01119_ clknet_leaf_278_clock u2.mem\[143\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10452_ _05029_ _05040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09444__I0 _04384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10980__S _05365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13171_ _01050_ clknet_leaf_264_clock u2.mem\[132\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10383_ _04993_ _00851_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06958__A1 u2.mem\[27\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12122_ _01485_ clknet_leaf_328_clock u2.select_mem_col\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_124_clock clknet_5_15_0_clock clknet_leaf_124_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_105_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12053_ net15 clknet_2_0__leaf_clock_a data_in_trans\[2\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06969__I _02447_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11004_ _05334_ _05380_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06186__A2 _01677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_139_clock clknet_5_13_0_clock clknet_leaf_139_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12955_ _00834_ clknet_leaf_198_clock u2.mem\[52\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11906_ _05945_ _01422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12886_ _00765_ clknet_leaf_63_clock u2.mem\[47\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07686__A2 _03088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11837_ _05876_ u2.mem\[189\]\[5\] _05895_ _05902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09683__I0 _04487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11768_ _05831_ u2.mem\[185\]\[2\] _05857_ _05860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11490__I0 _05677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13507_ _01386_ clknet_leaf_330_clock u2.mem\[188\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10719_ _05200_ u2.mem\[61\]\[2\] _05196_ _05201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11699_ _04120_ _05808_ _05817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11051__S _05403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08424__I _03753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13438_ _01317_ clknet_5_5_0_clock u2.mem\[176\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09435__I0 _04375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13369_ _01248_ clknet_leaf_356_clock u2.mem\[165\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_327_clock_I clknet_5_7_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09456__S _04419_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12429__CLK clknet_leaf_196_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07071__B1 _02549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07930_ u2.mem\[61\]\[14\] _02559_ _02561_ u2.mem\[63\]\[14\] _03395_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06879__I _02357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06964__A4 _02442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09255__I _04289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11545__I1 u2.mem\[171\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07861_ _02623_ _03328_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12579__CLK clknet_leaf_104_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07374__B2 u2.mem\[21\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09600_ _04509_ _00552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06812_ u2.mem\[179\]\[4\] _02151_ _02153_ u2.mem\[191\]\[4\] _02293_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07792_ _02460_ _03259_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09531_ _04118_ _04463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06743_ _02127_ _02226_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_3_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09462_ _04364_ u2.mem\[31\]\[3\] _04419_ _04423_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10130__S _04835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06674_ u2.mem\[146\]\[0\] _02156_ _02158_ u2.mem\[186\]\[0\] _02159_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08413_ _03672_ u2.mem\[7\]\[3\] _03754_ _03758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09393_ _04379_ _00475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11025__I _05394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08344_ _03710_ u2.mem\[5\]\[12\] _03711_ _03712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09674__I0 _04478_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10433__A1 _04180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08275_ _03491_ _03655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13204__CLK clknet_leaf_276_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07226_ u2.mem\[3\]\[2\] _02480_ _02359_ _02703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09426__I0 _04366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11896__S _05937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11233__I0 _05517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_41_clock clknet_5_6_0_clock clknet_leaf_41_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_164_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07157_ u2.mem\[45\]\[1\] _02633_ _02634_ u2.mem\[34\]\[1\] _02635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09366__S _04358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06108_ _01562_ _01574_ _01548_ _01615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_106_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13354__CLK clknet_leaf_359_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07088_ _02419_ _02567_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_65_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06039_ col_select_trans\[0\].data_sync col_select_trans\[1\].data_sync _01546_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10305__S _04944_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_56_clock clknet_5_12_0_clock clknet_leaf_56_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_87_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_51_clock_I clknet_5_13_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06168__A2 _01641_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09729_ _04589_ u2.mem\[37\]\[7\] _04580_ _04590_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10040__S _04777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12740_ _00619_ clknet_leaf_67_clock u2.mem\[38\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08509__I _03692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07413__I _02520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12671_ _00550_ clknet_leaf_177_clock u2.mem\[34\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_276_clock_I clknet_5_21_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11622_ _03487_ _05769_ _05770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09665__I0 _04469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11553_ _05717_ u2.mem\[171\]\[4\] _05721_ _05727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10504_ _05069_ _00896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09417__I0 _04356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11484_ _05668_ u2.mem\[167\]\[1\] _05683_ _05685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13223_ _01102_ clknet_leaf_286_clock u2.mem\[140\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10435_ _04987_ u2.mem\[54\]\[0\] _05030_ _05031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09276__S _04305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_7_0_clock clknet_0_clock clknet_3_7_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_174_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08180__S _03595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13154_ _01033_ clknet_leaf_263_clock u2.mem\[129\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10366_ _04913_ u2.mem\[52\]\[12\] _04981_ _04982_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08640__I1 u2.mem\[12\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12105_ _01488_ clknet_leaf_63_clock u2.active_mem\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10215__S _04887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13085_ _00964_ clknet_leaf_260_clock u2.mem\[60\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12721__CLK clknet_leaf_235_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10297_ _04920_ u2.mem\[50\]\[15\] _04938_ _04942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12036_ row_select_trans\[5\].A clknet_leaf_311_clock row_select_trans\[5\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06159__A2 _01665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07356__A1 _02821_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11152__A2 _05443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09803__I _04638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12871__CLK clknet_leaf_136_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10949__I _05345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07659__A2 _03049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06316__C1 u2.mem\[163\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12938_ _00817_ clknet_leaf_325_clock u2.mem\[50\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07323__I _02474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12088__D row_col_select_trans.A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12869_ _00748_ clknet_leaf_80_clock u2.mem\[46\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13227__CLK clknet_leaf_279_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09656__I0 _04498_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06390_ u2.mem\[175\]\[5\] _01601_ _01630_ u2.mem\[188\]\[5\] _01892_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_159_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08060_ _01945_ _03505_ _03514_ _00007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09408__I0 _04389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12251__CLK clknet_leaf_216_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07831__A2 _03139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07011_ u2.mem\[53\]\[0\] _02486_ _02489_ u2.mem\[56\]\[0\] _02490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11215__I0 _05514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11766__I1 u2.mem\[185\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09584__A2 _04441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08631__I1 u2.mem\[12\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08962_ _04019_ u2.mem\[20\]\[2\] _04097_ _04100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07913_ _03374_ _03375_ _03376_ _03377_ _03378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_64_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08893_ _04028_ u2.mem\[18\]\[6\] _04056_ _04059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07844_ _02592_ _03311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06555__C1 u2.mem\[181\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_9_0_clock clknet_4_4_0_clock clknet_5_9_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_84_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07775_ u2.mem\[6\]\[11\] _03094_ _03095_ u2.mem\[47\]\[11\] _03243_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09514_ _04375_ u2.mem\[32\]\[8\] _04453_ _04454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06726_ _02205_ _02206_ _02207_ _02208_ _02209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_52_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09445_ _04412_ _00494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06657_ _02141_ _02142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06322__A2 _01824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09376_ _04366_ u2.mem\[29\]\[4\] _04367_ _04368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09647__I0 _04489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_28_0_clock_I clknet_4_14_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06588_ u2.mem\[184\]\[0\] _02072_ _01994_ _02073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10257__I1 u2.mem\[49\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08327_ _03697_ _03698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07283__B1 _02667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08258_ _03563_ u2.mem\[4\]\[8\] _03645_ _03646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08064__I _03489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07209_ _02626_ _02687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08189_ _03577_ u2.mem\[2\]\[14\] _03600_ _03603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12744__CLK clknet_leaf_50_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10220_ _04575_ _04893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08622__I1 u2.mem\[12\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06389__A2 _01632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10151_ _04840_ _04851_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_79_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06794__C1 u2.mem\[159\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07408__I _02510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09824__S _04649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10082_ _04604_ _04810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12894__CLK clknet_leaf_214_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12124__CLK clknet_leaf_36_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08138__I0 _03570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06561__A2 _02036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08239__I _03634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10984_ _05346_ u2.mem\[136\]\[3\] _05365_ _05369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09886__I0 _04687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07143__I _02621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12723_ _00602_ clknet_leaf_71_clock u2.mem\[37\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11693__I0 _05794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12654_ _00533_ clknet_leaf_205_clock u2.mem\[33\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06982__I _02460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12274__CLK clknet_leaf_166_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09638__I0 _04480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11605_ _05759_ _01307_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12585_ _00464_ clknet_leaf_115_clock u2.mem\[28\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11536_ _05716_ _01281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07274__B1 _02489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07813__A2 _03123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11467_ _05672_ _01256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13206_ _01085_ clknet_leaf_271_clock u2.mem\[137\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10418_ _05018_ u2.mem\[53\]\[11\] _05012_ _05019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08702__I _03722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09810__I0 _04576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11398_ _05628_ _01231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07577__B2 u2.mem\[46\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13137_ _01016_ clknet_leaf_315_clock u2.mem\[63\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10349_ _04972_ _00838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07318__I _02460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09734__S _04593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06222__I _01565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13068_ _00947_ clknet_leaf_254_clock u2.mem\[59\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12019_ net31 clknet_2_2__leaf_clock_a mem_address_trans\[7\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09533__I _04464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07344__A4 _02818_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08129__I0 _03563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06552__A2 _02036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07560_ _02474_ _03031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12617__CLK clknet_leaf_111_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06511_ _01995_ _01996_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07491_ u2.mem\[5\]\[6\] _02920_ _02921_ u2.mem\[38\]\[6\] _02964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07501__A1 u2.mem\[27\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09230_ _04166_ _04278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06892__I _02370_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06442_ u2.mem\[194\]\[4\] _01924_ _01939_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09629__I0 _04471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09161_ _04232_ _00390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11436__I0 _05633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06373_ _01848_ _01853_ _01862_ _01875_ _01876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_33_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12767__CLK clknet_leaf_155_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08112_ _03552_ u2.mem\[1\]\[3\] _03546_ _03553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07002__B _02359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09092_ _04181_ _04192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_30_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07804__A2 _03114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08043_ _01769_ _03490_ _03501_ _00003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11739__I1 u2.mem\[183\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08612__I _03879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_224_clock_I clknet_5_25_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09994_ _04754_ _00701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06240__A1 u2.mem\[178\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06240__B2 u2.mem\[164\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08945_ _04073_ _04089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_83_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12147__CLK clknet_leaf_73_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06791__A2 _01995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08876_ _04048_ u2.mem\[17\]\[15\] _04042_ _04049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09443__I _04395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input22_I data_in_a[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07827_ _02553_ _03294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10589__I _03713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07758_ u2.mem\[60\]\[11\] _03055_ _03056_ u2.mem\[62\]\[11\] _03226_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12297__CLK clknet_leaf_120_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06709_ u2.mem\[180\]\[1\] _02043_ _02192_ u2.mem\[150\]\[1\] _02193_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13542__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07689_ _03155_ _03156_ _03157_ _03158_ _03159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_13_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09428_ _04369_ u2.mem\[30\]\[5\] _04401_ _04403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09359_ _04355_ _00465_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09245__A1 _04288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11213__I _03506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07256__B1 _02614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12370_ _00249_ clknet_leaf_150_clock u2.mem\[15\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11321_ _05552_ u2.mem\[157\]\[3\] _05576_ _05580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08522__I _03709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11252_ _05500_ u2.mem\[153\]\[0\] _05537_ _05538_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07559__B2 u2.mem\[7\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10203_ _04813_ u2.mem\[48\]\[13\] _04880_ _04882_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10402__I1 u2.mem\[53\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11183_ _05460_ u2.mem\[149\]\[0\] _05492_ _05493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07138__I _02616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06231__A1 u2.mem\[158\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10134_ _04782_ u2.mem\[47\]\[0\] _04841_ _04842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06231__B2 u2.mem\[151\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07574__A4 _03044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08359__I0 _03723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13072__CLK clknet_leaf_241_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10065_ _04798_ _00728_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06534__A2 _02018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07731__B2 u2.mem\[47\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10967_ _05343_ u2.mem\[135\]\[2\] _05356_ _05359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06298__A1 u2.mem\[146\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12706_ _00585_ clknet_leaf_238_clock u2.mem\[36\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10898_ _05313_ _01046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07601__I _02584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_173_clock_I clknet_5_27_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12637_ _00516_ clknet_leaf_192_clock u2.mem\[32\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07247__B1 _02587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12568_ _00447_ clknet_leaf_112_clock u2.mem\[27\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08633__S _03890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10962__I _05355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11519_ _05677_ u2.mem\[169\]\[4\] _05699_ _05705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12499_ _00378_ clknet_leaf_123_clock u2.mem\[23\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06470__A1 _01958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08598__I0 _03824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13415__CLK clknet_leaf_342_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07014__A3 _02392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06991_ _02466_ _02467_ _02468_ _02469_ _02470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11793__I _03679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06773__A2 _02252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08730_ _03955_ _00236_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07970__B2 u2.mem\[20\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06887__I _02365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_98_clock_I clknet_5_10_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08661_ _03910_ u2.mem\[13\]\[2\] _03906_ _03911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13565__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07612_ _02605_ _03083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08592_ _03817_ u2.mem\[11\]\[8\] _03867_ _03868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07543_ u2.mem\[45\]\[8\] _02866_ _02867_ u2.mem\[34\]\[8\] _03014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06289__A1 u2.mem\[190\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07486__B1 _02914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06289__B2 u2.mem\[194\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07474_ _02943_ _02944_ _02945_ _02946_ _02947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_39_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09213_ _04266_ _00408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11409__I0 _05635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06425_ _01545_ _01915_ _01921_ _01925_ _01458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09144_ _04221_ _00384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06356_ u2.mem\[159\]\[4\] _01603_ _01594_ u2.mem\[149\]\[4\] _01859_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08543__S _03836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07789__A1 u2.mem\[27\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09075_ _04119_ u2.mem\[22\]\[0\] _04182_ _04183_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06287_ u2.mem\[193\]\[2\] _01731_ _01734_ u2.mem\[177\]\[2\] _01792_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08026_ _03486_ _03487_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_146_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08342__I _03709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08589__I0 _03815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07005__A3 _02382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09977_ _04739_ _04745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_104_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11409__S _05624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08928_ _04023_ u2.mem\[19\]\[4\] _04079_ _04080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08859_ _03701_ _04037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07713__A1 u2.mem\[61\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_6_0_clock clknet_3_3_0_clock clknet_4_6_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_3658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11870_ _05923_ _01408_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08718__S _03947_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09901__I _04588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10821_ _05264_ _01018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11648__I0 _05758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11144__S _05462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10752_ _05222_ u2.mem\[61\]\[12\] _05223_ _05224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13540_ _01419_ clknet_leaf_34_clock u2.mem\[192\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13471_ _01350_ clknet_leaf_293_clock u2.mem\[182\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10683_ _05173_ _05179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_71_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12422_ _00301_ clknet_leaf_87_clock u2.mem\[18\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07229__B1 _02649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08453__S _03778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08816__I1 u2.mem\[16\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12353_ _00232_ clknet_leaf_150_clock u2.mem\[14\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10782__I _05231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12312__CLK clknet_leaf_121_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13438__CLK clknet_5_5_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11304_ _05570_ _01195_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12284_ _00163_ clknet_leaf_185_clock u2.mem\[10\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11235_ _05442_ _05527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_4_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09241__I1 u2.mem\[25\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06204__A1 u2.mem\[153\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06204__B2 u2.mem\[160\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11166_ _05442_ _05482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_121_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11319__S _05576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06755__A2 _02231_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10117_ _04804_ u2.mem\[46\]\[9\] _04830_ _04832_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11097_ _05439_ _01119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09083__I _04181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10048_ _04786_ u2.mem\[45\]\[1\] _04784_ _04787_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11887__I0 u2.mem\[192\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06507__A2 row_select_trans\[4\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08628__S _03885_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10957__I _05351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08504__I0 _03813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11999_ _00011_ clknet_leaf_28_clock u2.mem\[0\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07331__I _02485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10893__S _05310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06140__C2 _01646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06210_ _01706_ _01711_ _01716_ _01717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_129_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06691__B2 u2.mem\[161\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07190_ u2.mem\[61\]\[1\] _02666_ _02667_ u2.mem\[63\]\[1\] _02668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_157_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06141_ _01606_ _01628_ _01637_ _01647_ _01648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10692__I _05173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09480__I1 u2.mem\[31\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06443__A1 u2.mem\[193\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06072_ _01551_ _01579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06443__B2 u2.mem\[192\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09900_ _04697_ _00664_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10378__I0 _04987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08196__A1 _03605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09831_ _04605_ u2.mem\[39\]\[12\] _04654_ _04655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06746__A2 _02128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08991__I0 _04048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11229__S _05520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12955__CLK clknet_leaf_198_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09762_ _04614_ _04615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06974_ _02441_ _02421_ _02424_ _02453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XTAP_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07506__I _02358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08713_ _03912_ u2.mem\[14\]\[3\] _03942_ _03946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09693_ _04562_ _00592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11878__I0 u2.mem\[192\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08644_ _03831_ u2.mem\[12\]\[14\] _03895_ _03898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08575_ _03858_ _00178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09299__I1 u2.mem\[27\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07526_ u2.mem\[29\]\[7\] _02833_ _02834_ u2.mem\[11\]\[7\] _02998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08337__I _03705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07457_ u2.mem\[40\]\[6\] _02785_ _02786_ u2.mem\[30\]\[6\] _02930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12335__CLK clknet_leaf_152_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09369__S _04358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06682__A1 u2.mem\[185\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06408_ _01882_ _01887_ _01896_ _01909_ _01910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_155_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07388_ u2.mem\[6\]\[4\] _02861_ _02862_ u2.mem\[47\]\[4\] _02863_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06682__B2 u2.mem\[173\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11558__A2 _05729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09127_ _04151_ u2.mem\[23\]\[7\] _04208_ _04212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11802__I0 _05870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06339_ _01809_ _01555_ _01842_ _01483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09168__I _04225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09058_ _04169_ _00350_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12485__CLK clknet_leaf_100_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07631__B1 _03100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08072__I data_in_trans\[10\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07777__A4 _03244_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08009_ u2.active_mem\[3\] _03461_ _03462_ u2.active_mem\[2\] _03472_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_85_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11020_ _05391_ _01090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_121_clock_I clknet_5_15_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07529__A4 _03000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07934__A1 _03395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08982__I0 _04039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07416__I _02525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11869__I0 _05913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10978__S _05365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12971_ _00850_ clknet_leaf_246_clock u2.mem\[53\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08734__I0 _03932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07698__B1 _03029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11922_ _05954_ _01429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10541__I0 _05025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09631__I _04521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07162__A2 _02457_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11853_ _03674_ _05913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10804_ u2.mem\[63\]\[1\] _03497_ _05253_ _05255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11784_ _03666_ _05870_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_354_clock clknet_5_1_0_clock clknet_leaf_354_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_57_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13523_ _01402_ clknet_leaf_15_clock u2.mem\[190\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10735_ _05211_ u2.mem\[61\]\[7\] _05205_ _05212_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13260__CLK clknet_leaf_295_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_46_clock_I clknet_5_7_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06990__I _02362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10666_ _05124_ u2.mem\[59\]\[13\] _05167_ _05169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13454_ _01333_ clknet_leaf_300_clock u2.mem\[179\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12405_ _00284_ clknet_leaf_88_clock u2.mem\[17\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10218__S _04887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13385_ _01264_ clknet_leaf_306_clock u2.mem\[167\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10597_ _05129_ _00929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09462__I1 u2.mem\[31\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06425__A1 _01545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07100__B _02552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12336_ _00215_ clknet_leaf_222_clock u2.mem\[13\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07622__B1 _03092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08911__S _04066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12267_ _00146_ clknet_leaf_184_clock u2.mem\[9\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11218_ _05516_ _05517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12198_ _00077_ clknet_leaf_73_clock u2.mem\[4\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07925__A1 u2.mem\[14\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06728__A2 _02030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11049__S _05403_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08973__I0 _04030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07925__B2 u2.mem\[12\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11149_ _05351_ _05472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12208__CLK clknet_leaf_231_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10780__I0 _05211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07326__I _02479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09742__S _04593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_307_clock clknet_5_16_0_clock clknet_leaf_307_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_48_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08725__I0 _03923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06690_ _02107_ _02174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10532__I0 _05016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07153__A2 _02589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_323_clock_I clknet_5_18_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12358__CLK clknet_leaf_80_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08360_ _03724_ _00097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08157__I _03584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07061__I _02539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07311_ _02414_ _02786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08291_ _03668_ u2.mem\[5\]\[2\] _03660_ _03669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10835__I1 _05229_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08653__A2 _03904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06259__A4 _01764_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06664__A1 u2.mem\[170\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07242_ u2.mem\[57\]\[2\] _02554_ _02556_ u2.mem\[41\]\[2\] _02719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06664__B2 u2.mem\[156\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07173_ u2.mem\[53\]\[1\] _02486_ _02489_ u2.mem\[56\]\[1\] _02651_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10128__S _04835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08405__A2 _03752_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06124_ _01630_ _01631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06055_ col_select_trans\[0\].data_sync _01562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_132_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09716__I _04566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08964__I0 _04021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09814_ _04645_ _00630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10771__I0 _05202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06195__A3 _01580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13133__CLK clknet_leaf_268_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09745_ _04601_ _04602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06957_ _02435_ _02436_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08716__I0 _03914_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09676_ _04480_ u2.mem\[36\]\[7\] _04549_ _04553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06888_ _02339_ _02338_ _02344_ _02367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_54_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10523__I0 _05007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08627_ _03888_ _00200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13283__CLK clknet_leaf_360_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06352__C2 u2.mem\[168\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08558_ _03848_ _00171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09141__I0 _04171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07509_ u2.mem\[50\]\[7\] _02878_ _02879_ u2.mem\[51\]\[7\] _02981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_11_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10826__I1 _03525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08489_ _03803_ _00147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09099__S _04192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06655__A1 u2.mem\[154\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10520_ _05079_ _00902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06655__B2 u2.mem\[162\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10451_ _05039_ _00873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10038__S _04777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09444__I1 u2.mem\[30\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06407__A1 _01901_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13170_ _01049_ clknet_leaf_268_clock u2.mem\[131\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10382_ _04992_ u2.mem\[53\]\[1\] _04989_ _04993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06958__A2 _02428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12121_ _01484_ clknet_leaf_328_clock u2.select_mem_col\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12052_ data_in_trans\[1\].A clknet_leaf_287_clock data_in_trans\[1\].data_sync vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_272_clock_I clknet_5_20_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07907__A1 _03357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11003_ _05379_ _01085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06186__A3 _01580_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06050__I _01556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11891__I _05928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08707__I0 _03900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12500__CLK clknet_leaf_105_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10501__S _05066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08178__S _03595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10514__I0 _04995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12954_ _00833_ clknet_leaf_324_clock u2.mem\[51\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11905_ u2.mem\[192\]\[12\] _03528_ _05942_ _05945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_3_0_clock clknet_0_clock clknet_3_3_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_2540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12885_ _00764_ clknet_leaf_63_clock u2.mem\[47\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06343__C2 u2.mem\[181\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_293_clock clknet_5_20_0_clock clknet_leaf_293_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06894__A1 _02365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10300__I _04943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11836_ _05901_ _01396_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09132__I0 _04158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12650__CLK clknet_leaf_110_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10817__I1 _03515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11767_ _05859_ _01369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09683__I1 u2.mem\[36\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13506_ _01385_ clknet_leaf_330_clock u2.mem\[187\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10718_ _04994_ _05200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11698_ _05816_ _01343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13437_ _01316_ clknet_leaf_350_clock u2.mem\[176\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13006__CLK clknet_leaf_259_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10649_ _05159_ _00951_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09435__I1 u2.mem\[30\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11242__I1 u2.mem\[152\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06225__I _01577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13368_ _01247_ clknet_leaf_359_clock u2.mem\[164\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_231_clock clknet_5_24_0_clock clknet_leaf_231_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_6_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12319_ _00198_ clknet_leaf_157_clock u2.mem\[12\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13299_ _01178_ clknet_leaf_363_clock u2.mem\[153\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09199__I0 _04256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09536__I _04127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12030__CLK clknet_leaf_307_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08946__I0 _04041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07860_ _02621_ _03327_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_246_clock clknet_5_22_0_clock clknet_leaf_246_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_3_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06811_ u2.mem\[170\]\[4\] _02146_ _02148_ u2.mem\[156\]\[4\] _02292_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07791_ _02456_ _03258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12180__CLK clknet_leaf_75_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11507__S _05691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09530_ _04462_ _00529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06742_ _02126_ _02225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06895__I _02373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10505__I0 _05027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09461_ _04422_ _00500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06673_ _02157_ _02158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08412_ _03757_ _00116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09392_ _04378_ u2.mem\[29\]\[9\] _04376_ _04379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09123__I0 _04145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08343_ _03659_ _03711_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_33_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10808__I1 _03503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11242__S _05529_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08274_ _03654_ _00081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10433__A2 _04964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07225_ u2.mem\[16\]\[2\] _02475_ _02477_ u2.mem\[33\]\[2\] _02702_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_5_0_clock clknet_4_2_0_clock clknet_5_5_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_164_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09426__I1 u2.mem\[30\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09647__S _04532_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07156_ _02447_ _02634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11233__I1 u2.mem\[151\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06107_ _01567_ _01612_ _01613_ _01614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_105_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07062__A1 _02426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07087_ _02417_ _02566_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_161_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10992__I0 _05335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06038_ _01544_ _01545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_156_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08937__I0 _04032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12523__CLK clknet_leaf_183_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07989_ u2.mem\[39\]\[15\] _03321_ _03322_ u2.mem\[48\]\[15\] _03453_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11417__S _05638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09728_ _04588_ _04589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10321__S _04954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12673__CLK clknet_leaf_154_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09659_ _04095_ _04542_ _04543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_3_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06876__A1 _02339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12670_ _00549_ clknet_leaf_194_clock u2.mem\[34\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_219_clock_I clknet_5_28_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09114__I0 _04128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11621_ _05768_ _05769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13029__CLK clknet_leaf_31_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09665__I1 u2.mem\[36\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11552_ _05726_ _01287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10503_ _05025_ u2.mem\[55\]\[14\] _05066_ _05069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11483_ _05684_ _01260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12053__CLK clknet_2_0__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13222_ _01101_ clknet_leaf_280_clock u2.mem\[140\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13179__CLK clknet_leaf_275_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10434_ _05029_ _05030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_152_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07053__A1 _02454_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10365_ _04965_ _04981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_124_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13153_ _01032_ clknet_leaf_268_clock u2.mem\[129\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12104_ _01487_ clknet_leaf_63_clock u2.active_mem\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06800__A1 _02278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13084_ _00963_ clknet_leaf_261_clock u2.mem\[60\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10296_ _04941_ _00816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08928__I0 _04023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12035_ net42 clknet_2_3__leaf_clock_a row_select_trans\[5\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08002__B1 _03462_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10735__I0 _05211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09292__S _04313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06159__A3 _01591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_2_0_clock_I clknet_4_1_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07356__A2 _02824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10231__S _04896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12937_ _00816_ clknet_leaf_323_clock u2.mem\[50\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06316__B1 _01646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11160__I0 _05468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06316__C2 _01642_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06867__A1 _02338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12868_ _00747_ clknet_leaf_83_clock u2.mem\[46\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11819_ _05872_ u2.mem\[188\]\[3\] _05888_ _05892_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12799_ _00678_ clknet_leaf_144_clock u2.mem\[42\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11062__S _05413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07010_ _02488_ _02489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_170_clock clknet_5_27_0_clock clknet_leaf_170_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_31_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11215__I1 u2.mem\[150\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08371__S _03728_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12546__CLK clknet_leaf_168_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08961_ _04099_ _00323_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_185_clock clknet_5_30_0_clock clknet_leaf_185_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08919__I0 _04010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07912_ u2.mem\[27\]\[14\] _03254_ _03255_ u2.mem\[35\]\[14\] _03377_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08892_ _04058_ _00295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10726__I0 _05204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_168_clock_I clknet_5_27_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12696__CLK clknet_leaf_129_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09592__I0 _04471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07843_ _02590_ _03310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07774_ u2.mem\[8\]\[11\] _03091_ _03092_ u2.mem\[4\]\[11\] _03242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09513_ _04442_ _04453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06725_ u2.mem\[184\]\[2\] _02072_ _01995_ _02208_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06858__A1 _01878_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09444_ _04384_ u2.mem\[30\]\[12\] _04411_ _04412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06656_ _02064_ _02119_ _02141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_220_clock_I clknet_5_28_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_123_clock clknet_5_15_0_clock clknet_leaf_123_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09375_ _04357_ _04367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06587_ _02071_ _02072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12076__CLK clknet_leaf_343_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08326_ _03696_ _03697_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_28_0_clock clknet_4_14_0_clock clknet_5_28_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_20_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06293__C _01797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13321__CLK clknet_leaf_303_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08257_ _03634_ _03645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_21_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_138_clock clknet_5_13_0_clock clknet_leaf_138_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_20_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07208_ _02682_ _02683_ _02684_ _02685_ _02686_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_105_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08188_ _03602_ _00047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08281__S _03660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07139_ _02473_ _02438_ _02439_ _02384_ _02618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__10316__S _04949_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10965__I0 _05340_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07586__A2 _03055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10150_ _04850_ _00761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08080__I _03493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06794__B1 _02098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06794__C2 _02174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10081_ _04809_ _00733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07338__A2 _02654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11147__S _05461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10051__S _04784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10986__S _05364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10983_ _05368_ _01076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09886__I1 u2.mem\[41\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12722_ _00601_ clknet_leaf_235_clock u2.mem\[37\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08456__S _03783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06849__B2 u2.mem\[162\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12419__CLK clknet_leaf_110_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11693__I1 u2.mem\[180\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07510__A2 _02881_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12653_ _00532_ clknet_leaf_205_clock u2.mem\[33\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11604_ _05758_ u2.mem\[174\]\[5\] _05747_ _05759_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12584_ _00463_ clknet_leaf_115_clock u2.mem\[28\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07274__A1 u2.mem\[53\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12569__CLK clknet_leaf_113_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11535_ _05715_ u2.mem\[170\]\[3\] _05709_ _05716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07274__B2 u2.mem\[56\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11610__S _05761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08191__S _03600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11466_ _05671_ u2.mem\[166\]\[2\] _05665_ _05672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13205_ _01084_ clknet_leaf_275_clock u2.mem\[137\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10417_ _03704_ _05018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11397_ _05627_ u2.mem\[162\]\[1\] _05625_ _05628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07577__A2 _02893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13136_ _01015_ clknet_leaf_315_clock u2.mem\[63\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10348_ _04895_ u2.mem\[52\]\[4\] _04971_ _04972_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07041__A4 _02519_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10279_ _04902_ u2.mem\[50\]\[7\] _04928_ _04932_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13067_ _00946_ clknet_leaf_248_clock u2.mem\[59\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10708__I0 _05128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07329__A2 _02645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12018_ mem_address_trans\[6\].A clknet_leaf_299_clock mem_address_trans\[6\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11381__I0 _05587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07334__I _02494_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_40_clock clknet_5_6_0_clock clknet_leaf_40_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06510_ _01994_ _01995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07490_ _02959_ _02960_ _02961_ _02962_ _02963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_61_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06441_ _01914_ _01938_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09160_ _04140_ u2.mem\[24\]\[4\] _04231_ _04232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_55_clock clknet_5_12_0_clock clknet_leaf_55_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06372_ _01867_ _01868_ _01869_ _01874_ _01875_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__11436__I1 u2.mem\[164\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08111_ _03503_ _03552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_159_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09091_ _04191_ _00361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_94_clock_I clknet_5_10_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13494__CLK clknet_leaf_295_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08042_ _03500_ _03494_ _03501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10136__S _04841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06413__I _01913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09993_ _04707_ u2.mem\[43\]\[11\] _04750_ _04754_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06776__B1 _02078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08944_ _04088_ _00317_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08875_ _03722_ _04048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07826_ u2.mem\[37\]\[12\] _03291_ _03292_ u2.mem\[59\]\[12\] _03293_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_79_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09317__I0 _04283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input15_I data_in_a[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07757_ u2.mem\[61\]\[11\] _03132_ _03133_ u2.mem\[63\]\[11\] _03225_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11124__I0 _05426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06708_ _02047_ _02192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07688_ u2.mem\[6\]\[9\] _03094_ _03095_ u2.mem\[47\]\[9\] _03158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_77_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09427_ _04402_ _00486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06639_ u2.mem\[185\]\[0\] _02121_ _02123_ u2.mem\[173\]\[0\] _02124_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06700__B1 _02067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08075__I data_in_trans\[11\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09358_ _04285_ u2.mem\[28\]\[15\] _04351_ _04355_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09245__A2 _04250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08309_ data_in_trans\[6\].data_sync _03683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09289_ _04315_ _00435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11320_ _05579_ _01202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_2_0_clock clknet_3_1_0_clock clknet_4_2_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_165_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11251_ _05536_ _05537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_49_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10938__I0 _05335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07419__I _02530_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07559__A2 _03028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10202_ _04881_ _00782_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09835__S _04654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11182_ _05491_ _05492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_171_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07023__A4 _02393_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10133_ _04840_ _04841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__13217__CLK clknet_leaf_286_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09556__I0 _04480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10064_ _04797_ u2.mem\[45\]\[6\] _04793_ _04798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07192__B1 _02542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09308__I0 _04274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12241__CLK clknet_leaf_227_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07731__A2 _03094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13367__CLK clknet_leaf_354_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10966_ _05358_ _01069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12705_ _00584_ clknet_leaf_238_clock u2.mem\[36\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10897_ _05301_ u2.mem\[131\]\[2\] _05310_ _05313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_116_clock_I clknet_5_14_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12636_ _00515_ clknet_leaf_192_clock u2.mem\[32\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07247__A1 u2.mem\[28\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07247__B2 u2.mem\[31\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12567_ _00446_ clknet_leaf_113_clock u2.mem\[27\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_10_0_clock_I clknet_4_5_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11518_ _05704_ _01275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12498_ _00377_ clknet_leaf_161_clock u2.mem\[23\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06470__A2 _01955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11449_ _05659_ _01251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13119_ _00998_ clknet_leaf_243_clock u2.mem\[62\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_06990_ _02362_ _02469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_98_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09547__I0 _04473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input7_I data_in_a[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08660_ _03667_ _03910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07611_ u2.mem\[52\]\[8\] _03080_ _03081_ u2.mem\[21\]\[8\] _03082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08591_ _03856_ _03867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_148_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11106__I0 _05420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12734__CLK clknet_leaf_252_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07999__I _01665_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11515__S _05700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07542_ _02360_ _03013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07473_ u2.mem\[43\]\[6\] _02816_ _02817_ u2.mem\[20\]\[6\] _02946_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11314__I _05575_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09212_ _04265_ u2.mem\[25\]\[6\] _04261_ _04266_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11409__I1 u2.mem\[162\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06424_ u2.mem\[194\]\[0\] _01924_ _01925_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12884__CLK clknet_leaf_63_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07238__A1 _02699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09143_ _04174_ u2.mem\[23\]\[14\] _04218_ _04221_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08286__I0 _03664_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06355_ u2.mem\[175\]\[4\] _01601_ _01630_ u2.mem\[188\]\[4\] _01858_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10093__I0 _04817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09719__I _04143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09074_ _04181_ _04182_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_147_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06286_ u2.mem\[158\]\[2\] _01565_ _01572_ u2.mem\[151\]\[2\] _01589_ u2.mem\[168\]\[2\]
+ _01791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_50_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08025_ _03481_ _03482_ _03485_ _03486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_162_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_318_clock_I clknet_5_18_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09976_ _04744_ _00693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07410__B2 u2.mem\[56\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08927_ _04073_ _04079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_29_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11345__I0 _05595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08858_ _04036_ _00283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11896__I1 _03518_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07713__A2 _03132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07809_ _02499_ _03276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08789_ _03908_ u2.mem\[16\]\[1\] _03990_ _03992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10820_ u2.mem\[63\]\[8\] _03518_ _05263_ _05264_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10751_ _05195_ _05223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_125_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13470_ _01349_ clknet_leaf_347_clock u2.mem\[181\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10682_ _05178_ _00965_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12421_ _00300_ clknet_leaf_87_clock u2.mem\[18\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10084__I0 _04810_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12352_ _00231_ clknet_leaf_148_clock u2.mem\[14\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11303_ _05548_ u2.mem\[156\]\[1\] _05568_ _05570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12283_ _00162_ clknet_leaf_184_clock u2.mem\[10\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12607__CLK clknet_leaf_173_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11234_ _05526_ _01169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11584__I0 _05719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06988__I _02389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11165_ _05481_ _01145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09529__I0 _04391_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07952__A2 _02444_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06755__A3 _02232_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10116_ _04831_ _00746_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11096_ _05428_ u2.mem\[143\]\[3\] _05435_ _05439_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_42_clock_I clknet_5_6_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11336__I0 _05589_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10047_ _04569_ _04786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12757__CLK clknet_leaf_70_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08909__S _04066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11887__I1 _03507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07704__A2 _03039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07612__I _02605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11998_ _00010_ clknet_leaf_28_clock u2.mem\[0\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08504__I1 u2.mem\[9\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07468__A1 u2.mem\[58\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10949_ _05345_ _05346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11134__I _05461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_267_clock_I clknet_5_22_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06140__A1 u2.mem\[145\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06140__B2 u2.mem\[163\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12619_ _00498_ clknet_leaf_186_clock u2.mem\[31\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12137__CLK clknet_leaf_38_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06691__A2 _02096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09539__I _04131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06140_ u2.mem\[145\]\[0\] _01640_ _01643_ u2.mem\[163\]\[0\] u2.mem\[165\]\[0\]
+ _01646_ _01647_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_160_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07640__A1 _03106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06071_ u2.mem\[158\]\[0\] _01565_ _01572_ u2.mem\[151\]\[0\] _01577_ u2.mem\[193\]\[0\]
+ _01578_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_126_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12287__CLK clknet_leaf_164_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10378__I1 u2.mem\[53\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08196__A2 _03606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09830_ _04638_ _04654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_140_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08440__I0 _03723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08991__I1 u2.mem\[20\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09761_ data_in_trans\[15\].data_sync _04614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06973_ _02408_ _02452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08712_ _03945_ _00228_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09692_ _04496_ u2.mem\[36\]\[14\] _04559_ _04562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11878__I1 _03492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08643_ _03897_ _00207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08574_ _03798_ u2.mem\[11\]\[0\] _03857_ _03858_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07525_ u2.mem\[26\]\[7\] _02906_ _02907_ u2.mem\[10\]\[7\] _02997_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07456_ u2.mem\[32\]\[6\] _02782_ _02783_ u2.mem\[2\]\[6\] _02929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06407_ _01901_ _01902_ _01903_ _01908_ _01909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__13062__CLK clknet_leaf_30_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07387_ _02623_ _02862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09126_ _04211_ _00376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08353__I _03718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06338_ _01814_ _01819_ _01828_ _01841_ _01842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__11802__I1 u2.mem\[187\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09057_ _04167_ u2.mem\[21\]\[12\] _04168_ _04169_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06269_ u2.mem\[178\]\[2\] _01772_ _01773_ u2.mem\[164\]\[2\] _01774_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08008_ _03469_ _03470_ _03471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09759__I0 _04612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11566__I0 _05715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08431__I0 _03706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08982__I1 u2.mem\[20\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09959_ _04709_ u2.mem\[42\]\[12\] _04734_ _04735_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10123__I _04819_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12970_ _00849_ clknet_leaf_124_clock u2.mem\[52\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11869__I1 u2.mem\[191\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08734__I1 u2.mem\[14\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11921_ _05911_ u2.mem\[193\]\[3\] _05950_ _05954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06757__B _02239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10541__I1 u2.mem\[56\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11852_ _05912_ _01401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07432__I _02572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10803_ _05254_ _01010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08498__I0 _03808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10994__S _05373_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11783_ _05869_ _01375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13405__CLK clknet_leaf_304_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13522_ _01401_ clknet_leaf_16_clock u2.mem\[190\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06048__I _01554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10734_ _03687_ _05211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13453_ _01332_ clknet_leaf_301_clock u2.mem\[179\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10665_ _05168_ _00958_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12404_ _00283_ clknet_leaf_107_clock u2.mem\[17\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09998__I0 _04712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13384_ _01263_ clknet_leaf_301_clock u2.mem\[167\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10596_ _05128_ u2.mem\[57\]\[15\] _05122_ _05129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12335_ _00214_ clknet_leaf_152_clock u2.mem\[13\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07622__A1 u2.mem\[8\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06425__A2 _01915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07100__C _02455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07622__B2 u2.mem\[4\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12266_ _00145_ clknet_leaf_55_clock u2.mem\[8\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11217_ _03510_ _05516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10234__S _04896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08422__I0 _03689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06189__A1 _01685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12197_ _00076_ clknet_leaf_72_clock u2.mem\[4\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07607__I _02592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07925__A2 _02526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08973__I1 u2.mem\[20\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06511__I _01995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11148_ _05471_ _01138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11309__I0 _05554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10033__I _04761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11079_ _05345_ _05428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08725__I1 u2.mem\[14\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09922__I0 _04712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07153__A3 _02610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07342__I _02516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07310_ _02405_ _02785_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08374__S _03733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08290_ _03667_ _03668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06113__A1 _01619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07241_ u2.mem\[37\]\[2\] _02540_ _02542_ u2.mem\[59\]\[2\] _02718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10409__S _05012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10048__I0 _04786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09989__I0 _04703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07172_ u2.mem\[54\]\[1\] _02648_ _02649_ u2.mem\[55\]\[1\] _02650_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06123_ _01581_ _01629_ _01630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08661__I0 _03910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12922__CLK clknet_leaf_126_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06054_ _01560_ _01561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_156_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08413__I0 _03672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09813_ _04579_ u2.mem\[39\]\[4\] _04644_ _04645_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06719__A3 _02201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08964__I1 u2.mem\[20\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06421__I _01911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10920__A1 _04121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09744_ data_in_trans\[11\].data_sync _04601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06956_ _02429_ _02431_ _02433_ _02434_ _02435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_100_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_1_0_clock clknet_4_0_0_clock clknet_5_1_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_39_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09675_ _04552_ _00584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06887_ _02365_ _02366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12302__CLK clknet_leaf_181_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13428__CLK clknet_leaf_350_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08626_ _03813_ u2.mem\[12\]\[6\] _03885_ _03888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08348__I _03714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06352__A1 u2.mem\[158\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06352__B2 u2.mem\[151\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08557_ _03820_ u2.mem\[10\]\[9\] _03846_ _03848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09141__I1 u2.mem\[23\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07508_ _02975_ _02976_ _02977_ _02979_ _02980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_51_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08488_ _03802_ u2.mem\[9\]\[1\] _03800_ _03803_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12452__CLK clknet_leaf_84_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07301__B1 _02624_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13578__CLK clknet_leaf_37_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07439_ _02595_ _02913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07852__A1 _03309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06655__A2 _02126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10319__S _04954_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08083__I data_in_trans\[13\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10450_ _05009_ u2.mem\[54\]\[7\] _05035_ _05039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09109_ _04201_ _00369_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10381_ _04991_ _04992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12120_ _01483_ clknet_leaf_333_clock u2.select_mem_col\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_215_clock_I clknet_5_28_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10054__S _04784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12051_ net14 clknet_2_0__leaf_clock_a data_in_trans\[1\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07368__B1 _02681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07907__A2 _03362_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_4_2_0_clock_I clknet_3_1_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11002_ _05352_ u2.mem\[137\]\[5\] _05372_ _05379_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12953_ _00832_ clknet_leaf_324_clock u2.mem\[51\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11711__I0 _05798_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10514__I1 u2.mem\[56\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11904_ _05944_ _01421_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12884_ _00763_ clknet_leaf_63_clock u2.mem\[47\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06343__A1 u2.mem\[174\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06343__B2 u2.mem\[155\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11835_ _05874_ u2.mem\[189\]\[4\] _05895_ _05901_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11766_ _05829_ u2.mem\[185\]\[1\] _05857_ _05859_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07438__A4 _02911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13505_ _01384_ clknet_leaf_318_clock u2.mem\[187\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10717_ _05199_ _00979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08891__I0 _04026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11412__I _05637_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11697_ _05798_ u2.mem\[180\]\[5\] _05809_ _05816_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12945__CLK clknet_leaf_233_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07111__B _02463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13436_ _01315_ clknet_leaf_350_clock u2.mem\[176\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10648_ _05106_ u2.mem\[59\]\[5\] _05157_ _05159_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13367_ _01246_ clknet_leaf_354_clock u2.mem\[164\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10579_ _03700_ _05117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10450__I0 _05009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12318_ _00197_ clknet_leaf_199_clock u2.mem\[12\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06803__C1 u2.mem\[145\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07071__A2 _02546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13298_ _01177_ clknet_leaf_2_clock u2.mem\[153\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09199__I1 u2.mem\[25\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12249_ _00128_ clknet_leaf_55_clock u2.mem\[7\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10899__S _05310_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12325__CLK clknet_leaf_85_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06810_ u2.mem\[146\]\[4\] _02156_ _02158_ u2.mem\[186\]\[4\] _02291_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_151_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07790_ _03247_ _03250_ _03253_ _03256_ _03257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_96_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08369__S _03728_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09552__I _04147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06741_ u2.mem\[144\]\[2\] _02115_ _02117_ u2.mem\[182\]\[2\] _02224_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09460_ _04362_ u2.mem\[31\]\[2\] _04419_ _04422_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06672_ _02125_ _01999_ _02157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06334__A1 u2.mem\[146\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12475__CLK clknet_leaf_182_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07072__I _02347_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06334__B2 u2.mem\[186\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08411_ _03668_ u2.mem\[7\]\[2\] _03754_ _03757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09391_ _04157_ _04378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08342_ _03709_ _03710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08087__A1 _03533_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07800__I _02479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_164_clock_I clknet_5_26_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07834__A1 u2.mem\[29\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08273_ _03579_ u2.mem\[4\]\[15\] _03650_ _03654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06637__A2 _02018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08882__I0 _04017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07224_ u2.mem\[1\]\[2\] _02465_ _02471_ u2.mem\[7\]\[2\] _02701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07155_ _02443_ _02633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09727__I data_in_trans\[7\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06106_ _01593_ _01613_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10441__I0 _04998_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07086_ _02564_ _02565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13100__CLK clknet_leaf_264_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06037_ u2.mem\[0\]\[0\] _01544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09663__S _04544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_353_clock clknet_5_1_0_clock clknet_leaf_353_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08011__A1 _03472_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_24_0_clock clknet_4_12_0_clock clknet_5_24_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_59_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13250__CLK clknet_leaf_285_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10602__S _05131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07988_ u2.mem\[5\]\[15\] _02627_ _02629_ u2.mem\[38\]\[15\] _03452_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07770__B1 _03084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_89_clock_I clknet_5_10_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12818__CLK clknet_leaf_147_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09727_ data_in_trans\[7\].data_sync _04588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06939_ _02417_ _02418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_55_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10401__I _03683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09658_ _04440_ _04542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08078__I _03489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06325__A1 u2.mem\[144\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06325__B2 u2.mem\[182\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08609_ _03631_ _03774_ _03877_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_76_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06876__A2 _02354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09589_ _04503_ _00547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12968__CLK clknet_leaf_124_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11620_ _04861_ _05274_ _05768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_145_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11551_ _05715_ u2.mem\[171\]\[3\] _05722_ _05726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08873__I0 _04046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10502_ _05068_ _00895_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11482_ _05663_ u2.mem\[167\]\[0\] _05683_ _05684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11992__CLK clknet_leaf_329_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_306_clock clknet_5_16_0_clock clknet_leaf_306_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13221_ _01100_ clknet_leaf_281_clock u2.mem\[140\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10433_ _04180_ _04964_ _05029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13152_ _01031_ clknet_leaf_245_clock u2.mem\[128\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10364_ _04980_ _00845_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12348__CLK clknet_leaf_202_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12103_ _01501_ clknet_leaf_62_clock u2.active_mem\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13083_ _00962_ clknet_leaf_267_clock u2.mem\[60\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10295_ _04918_ u2.mem\[50\]\[14\] _04938_ _04941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08928__I1 u2.mem\[19\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08002__A1 u2.active_mem\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12034_ row_select_trans\[4\].A clknet_leaf_289_clock row_select_trans\[4\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06061__I col_select_trans\[3\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08002__B2 u2.active_mem\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11608__S _05761_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06996__I _02474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10512__S _05073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08189__S _03600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12498__CLK clknet_leaf_161_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_5_6_0_clock_I clknet_4_3_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10499__I0 _05020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12936_ _00815_ clknet_leaf_324_clock u2.mem\[50\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06316__B2 u2.mem\[165\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11160__I1 u2.mem\[147\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12867_ _00746_ clknet_leaf_60_clock u2.mem\[46\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11818_ _05891_ _01388_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12798_ _00677_ clknet_leaf_220_clock u2.mem\[42\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07620__I _02611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11749_ _05848_ _05849_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_72_1569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13123__CLK clknet_leaf_21_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13419_ _01298_ clknet_leaf_297_clock u2.mem\[173\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08960_ _04017_ u2.mem\[20\]\[1\] _04097_ _04099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13273__CLK clknet_leaf_9_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07067__I _02545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07911_ u2.mem\[40\]\[14\] _03251_ _03252_ u2.mem\[30\]\[14\] _03376_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_151_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08891_ _04026_ u2.mem\[18\]\[5\] _04056_ _04058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10726__I1 u2.mem\[61\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07842_ u2.mem\[23\]\[12\] _03146_ _03147_ u2.mem\[22\]\[12\] _03309_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_90_clock_I clknet_5_8_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06555__A1 u2.mem\[155\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07752__B1 _03124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06555__B2 u2.mem\[174\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06839__C _02318_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07773_ u2.mem\[39\]\[11\] _03088_ _03089_ u2.mem\[48\]\[11\] _03241_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09512_ _04452_ _00521_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06724_ u2.mem\[171\]\[2\] _02066_ _02068_ u2.mem\[157\]\[2\] _02207_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06307__A1 u2.mem\[167\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06307__B2 u2.mem\[183\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09443_ _04395_ _04411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_64_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06655_ u2.mem\[154\]\[0\] _02126_ _02127_ u2.mem\[162\]\[0\] _02139_ _02140_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XPHY_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09374_ _04139_ _04366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06586_ _02015_ _02070_ _02071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08325_ data_in_trans\[9\].data_sync _03696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08256_ _03644_ _00073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07283__A2 _02666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07207_ u2.mem\[18\]\[1\] _02606_ _02608_ u2.mem\[19\]\[1\] _02685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08607__I0 _03833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08187_ _03575_ u2.mem\[2\]\[13\] _03600_ _03602_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07138_ _02616_ _02617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09280__I0 _04285_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_292_clock clknet_5_20_0_clock clknet_leaf_292_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07069_ _02547_ _02371_ _02375_ _02411_ _02548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__06794__B2 u2.mem\[161\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12640__CLK clknet_leaf_172_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10080_ _04808_ u2.mem\[45\]\[11\] _04802_ _04809_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08535__A2 _03726_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10332__S _04959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09192__I _04251_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12790__CLK clknet_leaf_71_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10982_ _05343_ u2.mem\[136\]\[2\] _05365_ _05368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12721_ _00600_ clknet_leaf_235_clock u2.mem\[37\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_230_clock clknet_5_24_0_clock clknet_leaf_230_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09099__I0 _04164_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12652_ _00531_ clknet_leaf_205_clock u2.mem\[33\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08536__I _03835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12020__CLK clknet_leaf_289_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13146__CLK clknet_leaf_38_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07440__I _02597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11603_ _05679_ _05758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12583_ _00462_ clknet_leaf_115_clock u2.mem\[28\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_245_clock clknet_5_22_0_clock clknet_leaf_245_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_129_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11534_ _05673_ _05715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07274__A2 _02486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12170__CLK clknet_leaf_109_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11465_ _05670_ _05671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13204_ _01083_ clknet_leaf_276_clock u2.mem\[137\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10405__I0 _05009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10416_ _05017_ _00860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09271__I0 _04276_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11396_ _05504_ _05627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06234__B1 _01689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13135_ _01014_ clknet_leaf_314_clock u2.mem\[63\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10347_ _04965_ _04971_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06785__A1 u2.mem\[179\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06785__B2 u2.mem\[191\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_112_clock_I clknet_5_14_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13066_ _00945_ clknet_leaf_325_clock u2.mem\[58\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10278_ _04931_ _00808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12017_ net30 clknet_2_2__leaf_clock_a mem_address_trans\[6\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11381__I1 u2.mem\[161\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11137__I _05339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09830__I _04638_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12919_ _00798_ clknet_leaf_125_clock u2.mem\[49\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06440_ _01809_ _01915_ _01936_ _01937_ _01467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08446__I _03777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07350__I _02539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08837__I0 _04021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06371_ u2.mem\[147\]\[4\] _01675_ _01679_ u2.mem\[169\]\[4\] _01873_ _01874_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_159_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12513__CLK clknet_leaf_162_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08110_ _03551_ _00020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_37_clock_I clknet_5_6_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09090_ _04151_ u2.mem\[22\]\[7\] _04187_ _04191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08041_ _03499_ _03500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11600__I _05676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09262__I0 _04267_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12663__CLK clknet_leaf_58_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09992_ _04753_ _00700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06776__A1 u2.mem\[165\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06776__B2 u2.mem\[163\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07973__B1 _02561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08943_ _04039_ u2.mem\[19\]\[11\] _04084_ _04088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13019__CLK clknet_leaf_249_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11248__S _05528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10152__S _04851_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08874_ _04047_ _00288_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06528__A1 _02007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07725__B1 _03081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07825_ _02541_ _03292_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09317__I1 u2.mem\[27\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07756_ _03207_ _03213_ _03218_ _03223_ _03224_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_56_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08557__S _03846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12043__CLK clknet_2_2__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09740__I data_in_trans\[10\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11124__I1 u2.mem\[145\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06707_ u2.mem\[155\]\[1\] _02030_ _02035_ u2.mem\[174\]\[1\] u2.mem\[181\]\[1\]
+ _02039_ _02191_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA_clkbuf_leaf_314_clock_I clknet_5_19_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07687_ u2.mem\[8\]\[9\] _03091_ _03092_ u2.mem\[4\]\[9\] _03157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09426_ _04366_ u2.mem\[30\]\[4\] _04401_ _04402_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06638_ _02122_ _02123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08356__I data_in_trans\[15\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06700__A1 u2.mem\[171\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06700__B2 u2.mem\[157\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09357_ _04354_ _00464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08828__I0 _04010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12193__CLK clknet_leaf_228_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06569_ _02052_ _02053_ _02054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11711__S _05817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08308_ _03682_ _00087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07256__A2 _02612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09288_ _04254_ u2.mem\[27\]\[1\] _04313_ _04315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06464__B1 _01943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08239_ _03634_ _03635_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_166_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11250_ _04248_ _05527_ _05536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06604__I _02088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09253__I0 _04258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10201_ _04810_ u2.mem\[48\]\[12\] _04880_ _04881_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11060__I0 _05386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11181_ _04120_ _05482_ _05491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_122_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06767__B2 u2.mem\[152\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10132_ _04417_ _04760_ _04840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_69_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10063_ _04585_ _04797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09851__S _04666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07192__A1 u2.mem\[37\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09308__I1 u2.mem\[27\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08467__S _03788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10965_ _05340_ u2.mem\[135\]\[1\] _05356_ _05358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12536__CLK clknet_leaf_116_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12704_ _00583_ clknet_leaf_238_clock u2.mem\[36\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08266__I _03634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10874__I0 _05294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10896_ _05312_ _01045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07170__I _02508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_184_clock clknet_5_27_0_clock clknet_leaf_184_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12635_ _00514_ clknet_leaf_194_clock u2.mem\[32\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07247__A2 _02585_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12566_ _00445_ clknet_leaf_94_clock u2.mem\[27\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12686__CLK clknet_leaf_193_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11517_ _05674_ u2.mem\[169\]\[3\] _05700_ _05704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06455__B1 _01948_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12497_ _00376_ clknet_leaf_163_clock u2.mem\[23\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_199_clock clknet_5_28_0_clock clknet_leaf_199_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_7_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11448_ _05631_ u2.mem\[165\]\[3\] _05655_ _05659_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_5_14_0_clock_I clknet_4_7_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11051__I0 _05392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11379_ _05583_ u2.mem\[161\]\[0\] _05616_ _05617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06758__A1 u2.mem\[159\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06758__B2 u2.mem\[149\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13118_ _00997_ clknet_leaf_266_clock u2.mem\[62\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_122_clock clknet_5_15_0_clock clknet_leaf_122_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_112_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_263_clock_I clknet_5_23_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_2_2__f_clock_a_I clknet_0_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13049_ _00928_ clknet_leaf_45_clock u2.mem\[57\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07707__B1 _03121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12066__CLK clknet_leaf_32_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13311__CLK clknet_leaf_347_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07610_ _02602_ _03081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_137_clock clknet_5_13_0_clock clknet_leaf_137_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08590_ _03866_ _00185_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06930__A1 _02352_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11106__I1 u2.mem\[144\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07541_ _01951_ _02780_ _02991_ _03012_ _01499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_62_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13461__CLK clknet_leaf_344_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07486__A2 _02913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07472_ u2.mem\[49\]\[6\] _02893_ _02894_ u2.mem\[46\]\[6\] _02945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07080__I _02558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09211_ _04147_ _04265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06423_ _01923_ _01924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09142_ _04220_ _00383_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07238__A2 _02704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06354_ u2.mem\[187\]\[4\] _01633_ _01636_ u2.mem\[192\]\[4\] _01857_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09483__I0 _04384_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08286__I1 u2.mem\[5\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09001__S _04124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09073_ _04180_ _04122_ _04181_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11290__I0 _05550_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06285_ u2.mem\[145\]\[2\] _01639_ _01643_ u2.mem\[163\]\[2\] u2.mem\[165\]\[2\]
+ _01645_ _01790_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_159_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06997__A1 _02429_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09936__S _04719_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08024_ _03483_ _03484_ _03485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09235__I0 _04281_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06749__A1 u2.mem\[185\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09975_ _04689_ u2.mem\[43\]\[3\] _04740_ _04744_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08926_ _04078_ _00309_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11345__I1 u2.mem\[158\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08857_ _04035_ u2.mem\[17\]\[9\] _04033_ _04036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12559__CLK clknet_leaf_170_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07174__B2 u2.mem\[36\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07808_ _02494_ _03275_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08788_ _03991_ _00258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07739_ _03203_ _03204_ _03205_ _03206_ _03207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_2948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10750_ _03708_ _05222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08086__I data_in_trans\[14\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09409_ _04390_ _00480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10681_ _05101_ u2.mem\[60\]\[3\] _05174_ _05178_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12420_ _00299_ clknet_leaf_108_clock u2.mem\[18\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07229__A2 _02648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09474__I0 _04375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12351_ _00230_ clknet_leaf_148_clock u2.mem\[14\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09846__S _04661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11302_ _05569_ _01194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12282_ _00161_ clknet_leaf_119_clock u2.mem\[9\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08750__S _03963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11233_ _05517_ u2.mem\[151\]\[5\] _05519_ _05526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07874__B _03211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12089__CLK clknet_2_0__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11733__A1 _05354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11164_ _05472_ u2.mem\[147\]\[5\] _05474_ _05481_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13334__CLK clknet_leaf_5_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10115_ _04801_ u2.mem\[46\]\[8\] _04830_ _04831_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11095_ _05438_ _01118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_54_clock clknet_5_12_0_clock clknet_leaf_54_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11336__I1 u2.mem\[158\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10046_ _04785_ _00722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13484__CLK clknet_leaf_290_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11616__S _05760_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_69_clock clknet_5_9_0_clock clknet_leaf_69_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_95_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11997_ _00009_ clknet_leaf_33_clock u2.mem\[0\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10847__I0 _05200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10948_ _04134_ _05345_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06509__I _01993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08925__S _04074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06676__B1 _02144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10879_ _04994_ _05301_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_1461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11351__S _05598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12618_ _00497_ clknet_leaf_111_clock u2.mem\[30\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08724__I _03941_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09465__I0 _04366_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12549_ _00428_ clknet_leaf_98_clock u2.mem\[26\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06070_ _01552_ _01576_ _01577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_0_clock_I clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09555__I _04150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08196__A3 _03483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09760_ _04613_ _00608_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06972_ _02407_ _02451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__12701__CLK clknet_leaf_257_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07075__I _02553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08711_ _03910_ u2.mem\[14\]\[2\] _03942_ _03945_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09691_ _04561_ _00591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11526__S _05709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08642_ _03829_ u2.mem\[12\]\[13\] _03895_ _03897_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08573_ _03856_ _03857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_148_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07524_ _02992_ _02993_ _02994_ _02995_ _02996_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06419__I _01913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07455_ u2.mem\[45\]\[6\] _02866_ _02867_ u2.mem\[34\]\[6\] _02928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_168_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13207__CLK clknet_leaf_287_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06406_ u2.mem\[147\]\[5\] _01675_ _01679_ u2.mem\[169\]\[5\] _01907_ _01908_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09456__I0 _04356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07386_ _02621_ _02861_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09125_ _04148_ u2.mem\[23\]\[6\] _04208_ _04211_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06337_ _01829_ _01834_ _01835_ _01840_ _01841_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_157_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07092__B1 _02570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09056_ _04123_ _04168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12231__CLK clknet_leaf_52_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06154__I _01660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07631__A2 _03099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13357__CLK clknet_leaf_356_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06268_ _01620_ _01773_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08007_ u2.active_mem\[15\] _03461_ _03462_ u2.active_mem\[14\] _03470_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_89_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06199_ u2.mem\[190\]\[0\] _01703_ _01705_ u2.mem\[194\]\[0\] _01706_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05993__I row_col_select_trans.data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07919__B1 _02505_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11566__I1 u2.mem\[172\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_2_0_clock_I clknet_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07395__A1 u2.mem\[32\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12381__CLK clknet_leaf_206_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10404__I _03687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07934__A3 _03397_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09958_ _04718_ _04734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_131_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_159_clock_I clknet_5_26_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08909_ _04044_ u2.mem\[18\]\[13\] _04066_ _04068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09889_ _04689_ u2.mem\[41\]\[3\] _04683_ _04690_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11436__S _05646_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11920_ _05953_ _01428_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07698__A2 _03028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11851_ _05911_ u2.mem\[190\]\[3\] _05905_ _05912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11235__I _05442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10802_ u2.mem\[63\]\[0\] _03492_ _05253_ _05254_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_211_clock_I clknet_5_29_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11782_ _05868_ u2.mem\[186\]\[1\] _05866_ _05869_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08498__I1 u2.mem\[9\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13521_ _01400_ clknet_leaf_16_clock u2.mem\[190\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10733_ _05210_ _00984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11171__S _05484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13452_ _01331_ clknet_leaf_342_clock u2.mem\[178\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10664_ _05121_ u2.mem\[59\]\[12\] _05167_ _05168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07870__A2 _03333_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_19_0_clock clknet_4_9_0_clock clknet_5_19_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_12403_ _00282_ clknet_leaf_108_clock u2.mem\[17\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13383_ _01262_ clknet_leaf_301_clock u2.mem\[167\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10595_ _03721_ _05128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12334_ _00213_ clknet_leaf_206_clock u2.mem\[13\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07083__B1 _02561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08480__S _03793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07622__A2 _03091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12265_ _00144_ clknet_leaf_54_clock u2.mem\[8\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12724__CLK clknet_leaf_72_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09375__I _04357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11216_ _05515_ _01162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12196_ _00075_ clknet_leaf_71_clock u2.mem\[4\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11147_ _05470_ u2.mem\[146\]\[4\] _05461_ _05471_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11309__I1 u2.mem\[156\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11078_ _05427_ _01112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06948__B _02425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10029_ _04705_ u2.mem\[44\]\[10\] _04772_ _04775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07689__A2 _03156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07623__I _02621_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07153__A4 _02631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12104__CLK clknet_leaf_63_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08655__S _03906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06113__A2 _01607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07240_ u2.mem\[60\]\[2\] _02546_ _02549_ u2.mem\[62\]\[2\] _02717_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12254__CLK clknet_leaf_216_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07171_ _02510_ _02649_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06122_ _01558_ _01559_ _01585_ _01629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06053_ _01558_ _01559_ _01560_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09285__I _04312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06702__I _02100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09610__I0 _04489_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07377__B2 u2.mem\[19\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10224__I _04886_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09812_ _04638_ _04644_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06719__A4 _02202_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_160_clock_I clknet_5_26_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06955_ _02401_ _02391_ _02424_ _02434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_09743_ _04600_ _00604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11256__S _05537_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06858__B _02337_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09674_ _04478_ u2.mem\[36\]\[6\] _04549_ _04552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06886_ _01988_ _01997_ _02365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08625_ _03887_ _00199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07144__A4 _02453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11055__I _05412_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08556_ _03847_ _00170_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07507_ u2.mem\[3\]\[7\] _02801_ _02978_ _02979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11484__I0 _05668_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08487_ _03663_ _03802_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07438_ _02908_ _02909_ _02910_ _02911_ _02912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08364__I _03727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_20_0_clock clknet_4_10_0_clock clknet_5_20_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_126_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_85_clock_I clknet_5_11_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07369_ _02590_ _02844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12747__CLK clknet_leaf_216_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09108_ _04177_ u2.mem\[22\]\[15\] _04197_ _04201_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10380_ _04126_ _04991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09039_ _04123_ _04155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_139_1539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09195__I _04127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12050_ data_in_trans\[0\].A clknet_leaf_288_clock data_in_trans\[0\].data_sync vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12897__CLK clknet_leaf_224_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06612__I _02096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09601__I0 _04480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11001_ _05378_ _01084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07907__A3 _03367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12127__CLK clknet_leaf_36_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_6_0_clock_I clknet_3_3_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12952_ _00831_ clknet_leaf_49_clock u2.mem\[51\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11711__I1 u2.mem\[181\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06487__C _01964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11903_ u2.mem\[192\]\[11\] _03525_ _05942_ _05944_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12883_ _00762_ clknet_leaf_64_clock u2.mem\[47\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07540__A1 _02996_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12277__CLK clknet_leaf_102_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_362_clock_I clknet_5_0_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06059__I _01556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11834_ _05900_ _01395_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13522__CLK clknet_leaf_16_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11765_ _05858_ _01368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13504_ _01383_ clknet_leaf_331_clock u2.mem\[187\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10716_ _05198_ u2.mem\[61\]\[1\] _05196_ _05199_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11696_ _05815_ _01342_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10309__I _04943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13435_ _01314_ clknet_leaf_350_clock u2.mem\[176\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10647_ _05158_ _00950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07111__C _02544_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13366_ _01245_ clknet_leaf_359_clock u2.mem\[164\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10578_ _05116_ _00923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12317_ _00196_ clknet_leaf_197_clock u2.mem\[12\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13297_ _01176_ clknet_leaf_363_clock u2.mem\[153\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07618__I _02618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12248_ _00127_ clknet_leaf_55_clock u2.mem\[7\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06522__I _02006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10044__I _04783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12179_ _00058_ clknet_leaf_76_clock u2.mem\[3\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06031__B2 _01516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06582__A2 _02018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13052__CLK clknet_leaf_259_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06740_ _02219_ _02220_ _02221_ _02222_ _02223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_37_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07353__I _02553_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06671_ _02155_ _02156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08410_ _03756_ _00115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11804__S _05879_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09390_ _04377_ _00474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08385__S _03738_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08341_ _03708_ _03709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11466__I0 _05671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09284__A1 _04311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_107_clock_I clknet_5_11_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06098__A1 u2.mem\[175\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07295__B1 _02603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08184__I _03584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08272_ _03653_ _00080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06098__B2 u2.mem\[159\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07223_ u2.mem\[15\]\[2\] _02457_ _02461_ u2.mem\[13\]\[2\] _02700_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07154_ _01544_ _02361_ _02536_ _02632_ _01486_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09831__I0 _04605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06105_ _01561_ _01612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_106_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07085_ _02451_ _02452_ _02442_ _02544_ _02564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_12_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06036_ u3.data u3.enable net44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08398__I0 _03723_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08011__A2 _03473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input38_I row_select_a[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07987_ _03447_ _03448_ _03449_ _03450_ _03451_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_47_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06573__A2 _02036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07770__B2 u2.mem\[19\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06938_ _02387_ _02417_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09726_ _04587_ _00600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09657_ _04541_ _00577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06869_ _01579_ _01985_ _02348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_16_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08570__I0 _03833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08608_ _03876_ _00193_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_09588_ _04467_ u2.mem\[34\]\[1\] _04501_ _04503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08539_ _03802_ u2.mem\[10\]\[1\] _03836_ _03838_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11550_ _05725_ _01286_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07286__B1 _02556_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06607__I _02091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10501_ _05023_ u2.mem\[55\]\[13\] _05066_ _05068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11481_ _05682_ _05683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_109_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09918__I _04682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13220_ _01099_ clknet_leaf_282_clock u2.mem\[140\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10432_ _05028_ _00865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08822__I _03656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09822__I0 _04592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07589__A1 u2.mem\[37\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13151_ _01030_ clknet_leaf_269_clock u2.mem\[128\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10363_ _04911_ u2.mem\[52\]\[11\] _04976_ _04980_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_309_clock_I clknet_5_16_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12102_ _01500_ clknet_leaf_62_clock u2.active_mem\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06261__A1 _01745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13082_ _00961_ clknet_leaf_42_clock u2.mem\[59\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10294_ _04940_ _00815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08389__I0 _03706_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13075__CLK clknet_leaf_25_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12033_ net41 clknet_2_3__leaf_clock_a row_select_trans\[4\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10196__I0 _04806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08002__A2 _03461_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06013__A1 _01516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07761__A1 _03225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06564__A2 _02040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09889__I0 _04689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12935_ _00814_ clknet_leaf_49_clock u2.mem\[50\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07513__A1 _02981_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06316__A2 _01734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08561__I0 _03824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11624__S _05771_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12912__CLK clknet_leaf_147_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12866_ _00745_ clknet_leaf_151_clock u2.mem\[46\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11448__I0 _05631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11817_ _05870_ u2.mem\[188\]\[2\] _05888_ _05891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12797_ _00676_ clknet_leaf_220_clock u2.mem\[42\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07277__B1 _02655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11748_ _04223_ _05847_ _05848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_109_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11679_ _05805_ _01335_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13418_ _01297_ clknet_leaf_299_clock u2.mem\[173\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09813__I0 _04579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13418__CLK clknet_leaf_299_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13349_ _01228_ clknet_leaf_10_clock u2.mem\[161\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07348__I _02548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07910_ u2.mem\[32\]\[14\] _03248_ _03249_ u2.mem\[2\]\[14\] _03375_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08890_ _04057_ _00294_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10187__I0 _04797_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07841_ _03298_ _03301_ _03304_ _03307_ _03308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__12442__CLK clknet_leaf_128_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13568__CLK clknet_leaf_15_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_33_clock_I clknet_5_3_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07752__A1 u2.mem\[14\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06555__A2 _02030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07752__B2 u2.mem\[12\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07772_ u2.mem\[5\]\[11\] _03153_ _03154_ u2.mem\[38\]\[11\] _03240_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09511_ _04373_ u2.mem\[32\]\[7\] _04448_ _04452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06723_ u2.mem\[167\]\[2\] _02060_ _02062_ u2.mem\[183\]\[2\] _02206_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_168_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11687__I0 _05786_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08552__I0 _03815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12592__CLK clknet_leaf_168_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09442_ _04410_ _00493_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06654_ _02132_ _02135_ _02138_ _02139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_168_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09373_ _04365_ _00469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06585_ _02027_ _02001_ _02070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_258_clock_I clknet_5_23_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08324_ _03695_ _00090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07268__B1 _02477_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08255_ _03561_ u2.mem\[4\]\[7\] _03640_ _03644_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07206_ u2.mem\[52\]\[1\] _02601_ _02603_ u2.mem\[21\]\[1\] _02684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08186_ _03601_ _00046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08607__I1 u2.mem\[11\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09804__I0 _04565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07137_ _02568_ _02371_ _02375_ _02468_ _02616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_88_1566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07035__A3 _02433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_310_clock_I clknet_5_17_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09674__S _04549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07068_ _02347_ _02547_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_134_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06794__A2 _02096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11709__S _05817_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06019_ _01515_ _01522_ _01527_ _01516_ _01528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10178__I0 _04788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09473__I _04418_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08535__A3 _03776_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08791__I0 _03910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12935__CLK clknet_leaf_49_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08089__I data_in_trans\[15\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11678__I0 _05794_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09709_ _04574_ _00596_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10981_ _05367_ _01075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08543__I0 _03806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11444__S _05655_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12720_ _00599_ clknet_leaf_236_clock u2.mem\[37\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10350__I0 _04898_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12651_ _00530_ clknet_leaf_207_clock u2.mem\[33\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11602_ _05757_ _01306_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12582_ _00461_ clknet_leaf_100_clock u2.mem\[28\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08753__S _03968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11533_ _05714_ _01280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11464_ _03499_ _05670_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10415_ _05016_ u2.mem\[53\]\[10\] _05012_ _05017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13203_ _01082_ clknet_leaf_280_clock u2.mem\[137\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11395_ _05626_ _01230_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07168__I _02504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06234__A1 u2.mem\[170\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10346_ _04970_ _00837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06234__B2 u2.mem\[156\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13134_ _01013_ clknet_leaf_268_clock u2.mem\[63\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13065_ _00944_ clknet_leaf_47_clock u2.mem\[58\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10277_ _04900_ u2.mem\[50\]\[6\] _04928_ _04931_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10523__S _05078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12016_ mem_address_trans\[5\].A clknet_leaf_294_clock mem_address_trans\[5\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11905__I1 _03528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07734__A1 _01962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07498__B1 _02867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12918_ _00797_ clknet_leaf_84_clock u2.mem\[49\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10341__I0 _04889_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12849_ _00728_ clknet_leaf_154_clock u2.mem\[45\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11153__I _05474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06370_ _01870_ _01871_ _01872_ _01873_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06247__I _01592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_352_clock clknet_5_1_0_clock clknet_leaf_352_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09558__I _04153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08040_ data_in_trans\[2\].data_sync _03499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_174_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12808__CLK clknet_leaf_139_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13390__CLK clknet_leaf_355_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09991_ _04705_ u2.mem\[43\]\[10\] _04750_ _04753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11529__S _05709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06776__A2 _02075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07973__B2 u2.mem\[63\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08942_ _04087_ _00316_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12958__CLK clknet_leaf_197_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07806__I _02488_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08873_ _04046_ u2.mem\[17\]\[14\] _04042_ _04047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06528__A2 _02012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08773__I0 _03935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07824_ _02539_ _03291_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10580__I0 _05117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07755_ _03219_ _03220_ _03221_ _03222_ _03223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xclkbuf_leaf_305_clock clknet_5_16_0_clock clknet_leaf_305_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_53_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06706_ _02184_ _02188_ _02189_ _02190_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07686_ u2.mem\[39\]\[9\] _03088_ _03089_ u2.mem\[48\]\[9\] _03156_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10332__I0 _04918_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09425_ _04395_ _04401_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_25_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06637_ _02064_ _02018_ _02122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12338__CLK clknet_leaf_152_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06700__A2 _02065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09356_ _04283_ u2.mem\[28\]\[14\] _04351_ _04354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06568_ _01998_ _02053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08307_ _03681_ u2.mem\[5\]\[5\] _03677_ _03682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09287_ _04314_ _00434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06499_ row_select_trans\[0\].data_sync _01984_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08238_ _03630_ _03542_ _03633_ _03634_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__06464__A1 u2.mem\[193\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12488__CLK clknet_leaf_164_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06464__B2 u2.mem\[194\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08169_ _03557_ u2.mem\[2\]\[5\] _03590_ _03592_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10407__I _03691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10399__I0 _05005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10200_ _04864_ _04880_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06216__A1 u2.mem\[173\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06216__B2 u2.mem\[185\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11180_ _05490_ _01151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07964__A1 u2.mem\[53\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10131_ _04839_ _00753_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10343__S _04966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10062_ _04796_ _00727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08764__I0 _03926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10142__I _04840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08748__S _03963_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09931__I _04718_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07192__A2 _02540_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13113__CLK clknet_leaf_327_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10323__I0 _04909_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10964_ _05357_ _01068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12703_ _00582_ clknet_leaf_239_clock u2.mem\[36\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07495__A3 _02966_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13263__CLK clknet_leaf_272_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10895_ _05299_ u2.mem\[131\]\[1\] _05310_ _05312_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12634_ _00513_ clknet_leaf_114_clock u2.mem\[31\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06067__I col_select_trans\[1\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11823__I0 _05876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12565_ _00444_ clknet_leaf_96_clock u2.mem\[27\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09378__I _04144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07652__B1 _03121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11516_ _05703_ _01274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12496_ _00375_ clknet_leaf_163_clock u2.mem\[23\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11447_ _05658_ _01250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11378_ _05615_ _05616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06758__A2 _02174_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_206_clock_I clknet_5_29_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11349__S _05598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10329_ _04960_ _00830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13117_ _00996_ clknet_leaf_261_clock u2.mem\[62\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_5_18_0_clock_I clknet_4_9_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13048_ _00927_ clknet_leaf_44_clock u2.mem\[57\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07707__A1 u2.mem\[44\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08755__I0 _03917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08658__S _03906_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09841__I _04660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08507__I0 _03815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06391__B1 _01594_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06930__A2 _02376_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07540_ _02996_ _03001_ _03006_ _03011_ _03012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_53_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10314__I0 _04900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07361__I _02579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09180__I0 _04171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07471_ u2.mem\[14\]\[6\] _02890_ _02891_ u2.mem\[12\]\[6\] _02944_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_291_clock clknet_5_20_0_clock clknet_leaf_291_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_62_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09210_ _04264_ _00407_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06422_ _01922_ _01916_ _01923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06694__A1 u2.mem\[149\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12630__CLK clknet_leaf_96_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09141_ _04171_ u2.mem\[23\]\[13\] _04218_ _04220_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06353_ u2.mem\[193\]\[4\] _01731_ _01734_ u2.mem\[177\]\[4\] _01856_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07238__A3 _02709_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09072_ _04179_ _04180_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_120_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07643__B1 _03112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11290__I1 u2.mem\[155\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06284_ u2.mem\[166\]\[2\] _01753_ _01754_ u2.mem\[161\]\[2\] _01788_ _01789_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_163_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06997__A2 _02445_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08023_ mem_write_n_trans.data_sync mem_address_trans\[9\].data_sync mem_address_trans\[8\].data_sync
+ _03484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_30_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10227__I _04582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12780__CLK clknet_leaf_253_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10163__S _04856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09974_ _04743_ _00692_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12010__CLK clknet_leaf_312_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09952__S _04729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08925_ _04021_ u2.mem\[19\]\[3\] _04074_ _04078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08746__I0 _03908_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08856_ _03697_ _04035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input20_I data_in_a[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_244_clock clknet_5_19_0_clock clknet_leaf_244_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07174__A2 _02495_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07807_ u2.mem\[53\]\[12\] _03272_ _03273_ u2.mem\[56\]\[12\] _03274_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_3639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12160__CLK clknet_leaf_152_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08787_ _03900_ u2.mem\[16\]\[0\] _03990_ _03991_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05999_ _01507_ _01508_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07738_ u2.mem\[27\]\[11\] _03021_ _03022_ u2.mem\[35\]\[11\] _03206_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10305__I0 _04891_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09171__I0 _04158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_259_clock clknet_5_23_0_clock clknet_leaf_259_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_164_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07669_ _02572_ _03139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09408_ _04389_ u2.mem\[29\]\[14\] _04385_ _04390_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07882__B1 _02528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10680_ _05177_ _00964_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_2_clock_I clknet_5_0_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_155_clock_I clknet_5_27_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09339_ _04344_ _00456_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09474__I1 u2.mem\[31\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09198__I _04131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06437__A1 _01769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07634__B1 _03022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12350_ _00229_ clknet_leaf_201_clock u2.mem\[14\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06437__B2 _01935_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11301_ _05544_ u2.mem\[156\]\[0\] _05568_ _05569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12281_ _00160_ clknet_leaf_119_clock u2.mem\[9\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11232_ _05525_ _01168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08830__I _03663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07937__A1 u2.mem\[9\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08985__I0 _04041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11733__A2 _05808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11169__S _05484_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11163_ _05480_ _01144_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10792__I0 _05222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07446__I _02626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09862__S _04671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10114_ _04819_ _04830_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_96_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11094_ _05426_ u2.mem\[143\]\[2\] _05435_ _05438_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12503__CLK clknet_leaf_121_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_15_0_clock clknet_4_7_0_clock clknet_5_15_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_10045_ _04782_ u2.mem\[45\]\[0\] _04784_ _04785_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08478__S _03793_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07165__A2 _02480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08277__I _03656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11996_ _00008_ clknet_leaf_320_clock u2.mem\[0\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09162__I0 _04145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12653__CLK clknet_leaf_205_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10947_ _05344_ _01064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11632__S _05770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06676__A1 u2.mem\[169\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06676__B2 u2.mem\[147\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10878_ _05300_ _01039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09102__S _04197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12617_ _00496_ clknet_leaf_111_clock u2.mem\[30\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13009__CLK clknet_leaf_239_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07625__B1 _03095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06525__I row_select_trans\[3\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12548_ _00427_ clknet_leaf_98_clock u2.mem\[26\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08941__S _04084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12479_ _00358_ clknet_leaf_163_clock u2.mem\[22\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12033__CLK clknet_2_3__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13159__CLK clknet_leaf_274_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08976__I0 _04032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_357_clock_I clknet_5_1_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10783__I0 _05213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06971_ _02397_ _02416_ _02437_ _02449_ _02450_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_98_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12183__CLK clknet_leaf_61_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08710_ _03944_ _00227_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09690_ _04494_ u2.mem\[36\]\[13\] _04559_ _04561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09571__I _04166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08641_ _03896_ _00206_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06364__B1 _01701_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08572_ _03605_ _03606_ _03607_ _03776_ _03856_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__07091__I _02569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09153__I0 _04128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07523_ u2.mem\[57\]\[7\] _02828_ _02829_ u2.mem\[41\]\[7\] _02995_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08900__I0 _04035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07454_ _01877_ _02780_ _02898_ _02927_ _01497_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06667__A1 _02104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06405_ _01904_ _01905_ _01906_ _01907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06863__C col_select_trans\[4\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10158__S _04851_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07385_ u2.mem\[8\]\[4\] _02858_ _02859_ u2.mem\[4\]\[4\] _02860_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_10_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09456__I1 u2.mem\[31\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11341__I _05513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09124_ _04210_ _00375_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07616__B1 _02921_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06336_ u2.mem\[147\]\[3\] _01676_ _01680_ u2.mem\[169\]\[3\] _01839_ _01840_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_148_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07092__A1 u2.mem\[29\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09055_ _04166_ _04167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06267_ _01618_ _01772_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08006_ u2.active_mem\[12\] _03458_ _03459_ u2.active_mem\[13\] _03469_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_102_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06198_ _01704_ _01705_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08967__I0 _04023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12526__CLK clknet_leaf_187_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10774__I0 _05204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09957_ _04733_ _00685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_183_clock clknet_5_30_0_clock clknet_leaf_183_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_4104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08908_ _04067_ _00302_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_6_0_clock_I clknet_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09888_ _04575_ _04689_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_81_clock_I clknet_5_8_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09392__I0 _04378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12676__CLK clknet_leaf_90_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08839_ _03675_ _04023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06355__B1 _01630_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10420__I _03708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11850_ _03670_ _05911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_166_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_198_clock clknet_5_30_0_clock clknet_leaf_198_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10801_ _05252_ _05253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_122_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10829__I1 _03528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11781_ _03662_ _05868_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11452__S _05654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06658__A1 _02023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13520_ _01399_ clknet_leaf_16_clock u2.mem\[190\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11651__A1 _05295_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10732_ _05209_ u2.mem\[61\]\[6\] _05205_ _05210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_121_clock clknet_5_15_0_clock clknet_leaf_121_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_15_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13451_ _01330_ clknet_leaf_342_clock u2.mem\[178\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10663_ _05151_ _05167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11251__I _05536_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12402_ _00281_ clknet_leaf_155_clock u2.mem\[17\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09857__S _04666_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11254__I1 u2.mem\[153\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13382_ _01261_ clknet_leaf_309_clock u2.mem\[167\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10594_ _05127_ _00928_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07083__A1 u2.mem\[61\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12333_ _00212_ clknet_leaf_209_clock u2.mem\[13\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_136_clock clknet_5_13_0_clock clknet_leaf_136_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_147_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06830__A1 u2.mem\[150\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12264_ _00143_ clknet_leaf_65_clock u2.mem\[8\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08958__I0 _04010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11215_ _05514_ u2.mem\[150\]\[4\] _05501_ _05515_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12195_ _00074_ clknet_leaf_72_clock u2.mem\[4\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13451__CLK clknet_leaf_342_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10765__I0 _05194_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07176__I _02520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09592__S _04501_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11146_ _05348_ _05470_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11077_ _05426_ u2.mem\[142\]\[2\] _05422_ _05427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09391__I _04157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06948__C _02426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10028_ _04774_ _00715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11979_ _05987_ _01453_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06649__A1 _01999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09767__S _04618_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07170_ _02508_ _02648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08671__S _03915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06121_ u2.mem\[171\]\[0\] _01611_ _01614_ u2.mem\[157\]\[0\] _01627_ _01628_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07074__A1 _02551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12549__CLK clknet_leaf_98_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06821__A1 u2.mem\[185\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06052_ col_select_trans\[3\].data_sync _01559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07086__I _02564_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09811_ _04643_ _00629_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_103_clock_I clknet_5_11_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09742_ _04599_ u2.mem\[37\]\[10\] _04593_ _04600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10441__S _05030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06954_ _02432_ _02433_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09673_ _04551_ _00583_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06885_ _02363_ _02364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_94_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08624_ _03811_ u2.mem\[12\]\[5\] _03885_ _03887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06888__A1 _02339_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08555_ _03817_ u2.mem\[10\]\[8\] _03846_ _03847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07506_ _02358_ _02978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12079__CLK clknet_2_1__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08486_ _03801_ _00146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11484__I1 u2.mem\[167\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13324__CLK clknet_leaf_342_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07301__A2 _02622_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07437_ u2.mem\[28\]\[5\] _02839_ _02840_ u2.mem\[31\]\[5\] _02911_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07852__A3 _03315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_13_0_clock_I clknet_3_6_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_28_clock_I clknet_5_3_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_53_clock clknet_5_12_0_clock clknet_leaf_53_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_13_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07368_ u2.mem\[23\]\[4\] _02680_ _02681_ u2.mem\[22\]\[4\] _02843_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09107_ _04200_ _00368_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06319_ u2.mem\[175\]\[3\] _01602_ _01631_ u2.mem\[188\]\[3\] _01823_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07299_ u2.mem\[39\]\[3\] _02617_ _02619_ u2.mem\[48\]\[3\] _02775_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06812__A1 u2.mem\[179\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09038_ _04153_ _04154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06812__B2 u2.mem\[191\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_68_clock clknet_5_9_0_clock clknet_leaf_68_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_85_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07368__A2 _02680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11000_ _05349_ u2.mem\[137\]\[4\] _05372_ _05378_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07907__A4 _03372_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12951_ _00830_ clknet_leaf_49_clock u2.mem\[51\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06328__B1 _01714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11902_ _05943_ _01420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12882_ _00761_ clknet_leaf_230_clock u2.mem\[47\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07540__A2 _03001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_305_clock_I clknet_5_16_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11833_ _05872_ u2.mem\[189\]\[3\] _05896_ _05900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11764_ _05825_ u2.mem\[185\]\[0\] _05857_ _05858_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13503_ _01382_ clknet_leaf_331_clock u2.mem\[187\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10715_ _04991_ _05198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11695_ _05796_ u2.mem\[180\]\[4\] _05809_ _05815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11227__I1 u2.mem\[151\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13434_ _01313_ clknet_leaf_337_clock u2.mem\[175\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08491__S _03800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10646_ _05103_ u2.mem\[59\]\[4\] _05157_ _05158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13365_ _01244_ clknet_leaf_358_clock u2.mem\[164\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10577_ _05115_ u2.mem\[57\]\[9\] _05113_ _05116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10986__I0 _05349_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12316_ _00195_ clknet_leaf_200_clock u2.mem\[12\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08290__I _03667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06803__A1 u2.mem\[165\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06803__B2 u2.mem\[163\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13296_ _01175_ clknet_leaf_7_clock u2.mem\[152\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12247_ _00126_ clknet_leaf_55_clock u2.mem\[7\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12178_ _00057_ clknet_leaf_225_clock u2.mem\[3\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11357__S _05597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11129_ _05458_ _01132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12991__CLK clknet_leaf_239_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09356__I0 _04283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06319__B1 _01631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10060__I _04582_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06670_ _02108_ _02052_ _02155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12221__CLK clknet_leaf_213_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10910__I0 _05299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09108__I0 _04177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13347__CLK clknet_leaf_17_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11092__S _05435_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08340_ data_in_trans\[12\].data_sync _03708_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09284__A2 _04250_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07295__A1 u2.mem\[52\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08271_ _03577_ u2.mem\[4\]\[14\] _03650_ _03653_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12371__CLK clknet_leaf_78_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13497__CLK clknet_leaf_316_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07222_ _02695_ _02696_ _02697_ _02698_ _02699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_160_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07153_ _02563_ _02589_ _02610_ _02631_ _02632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_160_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07809__I _02499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06104_ _01610_ _01611_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07084_ _02543_ _02550_ _02557_ _02562_ _02563_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_156_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07062__A4 _02425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06035_ _01543_ _00000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10729__I0 _05207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09595__I0 _04473_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_254_clock_I clknet_5_23_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11267__S _05546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07986_ u2.mem\[18\]\[15\] _03316_ _03317_ u2.mem\[19\]\[15\] _03450_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_75_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07544__I _02385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09347__I0 _04274_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07770__A2 _03083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09725_ _04586_ u2.mem\[37\]\[6\] _04580_ _04587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06937_ u2.mem\[40\]\[0\] _02406_ _02415_ u2.mem\[30\]\[0\] _02416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11154__I0 _05460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09656_ _04498_ u2.mem\[35\]\[15\] _04537_ _04541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08576__S _03857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06868_ _02346_ _02347_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10901__I0 _05305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08570__I1 u2.mem\[10\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08607_ _03833_ u2.mem\[11\]\[15\] _03872_ _03876_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09587_ _04502_ _00546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_06799_ u2.mem\[184\]\[4\] _02071_ _01993_ _02280_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12714__CLK clknet_leaf_49_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05999__I _01507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08538_ _03837_ _00162_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11606__A1 _04416_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08469_ _03702_ u2.mem\[8\]\[10\] _03788_ _03791_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06628__A4 _02112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10500_ _05067_ _00894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11480_ _05354_ _05645_ _05682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__12864__CLK clknet_leaf_148_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10431_ _05027_ u2.mem\[53\]\[15\] _05021_ _05028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06623__I _02022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13150_ _01029_ clknet_leaf_262_clock u2.mem\[128\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10362_ _04979_ _00844_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07053__A4 _02411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12101_ _01499_ clknet_leaf_144_clock u2.active_mem\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06261__A2 _01751_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10293_ _04916_ u2.mem\[50\]\[13\] _04938_ _04940_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13081_ _00960_ clknet_leaf_40_clock u2.mem\[59\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09586__I0 _04463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12032_ row_select_trans\[3\].A clknet_leaf_302_clock row_select_trans\[3\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11177__S _05483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12244__CLK clknet_leaf_74_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09338__I0 _04265_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12012__D mem_address_trans\[3\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11905__S _05942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12934_ _00813_ clknet_leaf_31_clock u2.mem\[50\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12865_ _00744_ clknet_leaf_148_clock u2.mem\[46\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06721__B1 _02171_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08285__I _03663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11816_ _05890_ _01387_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11448__I1 u2.mem\[165\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12796_ _00675_ clknet_leaf_220_clock u2.mem\[42\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11747_ _05768_ _05847_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11640__S _05779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11678_ _05794_ u2.mem\[179\]\[3\] _05801_ _05805_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07029__A1 _02413_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13417_ _01296_ clknet_leaf_298_clock u2.mem\[173\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10629_ _05124_ u2.mem\[58\]\[13\] _05146_ _05148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07629__I _02443_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13348_ _01227_ clknet_leaf_17_clock u2.mem\[161\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06252__A2 _01755_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13279_ _01158_ clknet_leaf_361_clock u2.mem\[150\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07840_ u2.mem\[28\]\[12\] _03305_ _03306_ u2.mem\[31\]\[12\] _03307_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07364__I _02584_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09329__I0 _04256_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07752__A2 _03123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07771_ _03235_ _03236_ _03237_ _03238_ _03239_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_110_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09510_ _04451_ _00520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12737__CLK clknet_leaf_232_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11815__S _05888_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06722_ u2.mem\[164\]\[2\] _02051_ _02055_ u2.mem\[178\]\[2\] _02205_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11687__I1 u2.mem\[180\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08552__I1 u2.mem\[10\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09441_ _04382_ u2.mem\[30\]\[11\] _04406_ _04410_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06653_ u2.mem\[153\]\[0\] _02136_ _02137_ u2.mem\[160\]\[0\] _02138_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_91_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09372_ _04364_ u2.mem\[29\]\[3\] _04358_ _04365_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08195__I _03541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06708__I _02047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06584_ u2.mem\[171\]\[0\] _02066_ _02068_ u2.mem\[157\]\[0\] _02069_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12887__CLK clknet_leaf_57_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08323_ _03693_ u2.mem\[5\]\[8\] _03694_ _03695_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08254_ _03643_ _00072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07205_ u2.mem\[17\]\[1\] _02591_ _02593_ u2.mem\[24\]\[1\] _02683_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12117__CLK clknet_leaf_332_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06491__A2 _01917_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08185_ _03572_ u2.mem\[2\]\[12\] _03600_ _03601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07136_ u2.mem\[8\]\[0\] _02612_ _02614_ u2.mem\[4\]\[0\] _02615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07035__A4 _02425_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06779__B1 _02013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07067_ _02545_ _02546_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06018_ _01504_ _01524_ _01526_ _01527_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13512__CLK clknet_leaf_330_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11375__I0 _05595_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08240__I0 _03539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07969_ u2.mem\[49\]\[15\] _02531_ _02533_ u2.mem\[46\]\[15\] _03433_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09708_ _04573_ u2.mem\[37\]\[2\] _04567_ _04574_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11678__I1 u2.mem\[179\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10980_ _05340_ u2.mem\[136\]\[1\] _05365_ _05367_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09639_ _04531_ _00569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12650_ _00529_ clknet_leaf_110_clock u2.mem\[32\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07259__A1 _02720_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11601_ _05756_ u2.mem\[174\]\[4\] _05747_ _05757_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12581_ _00460_ clknet_leaf_98_clock u2.mem\[28\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11532_ _05713_ u2.mem\[170\]\[2\] _05709_ _05714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08833__I _03667_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11463_ _05669_ _01255_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13042__CLK clknet_leaf_321_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06482__A2 _01929_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13202_ _01081_ clknet_leaf_280_clock u2.mem\[137\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10414_ _03700_ _05016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11394_ _05623_ u2.mem\[162\]\[0\] _05625_ _05626_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13133_ _01012_ clknet_leaf_268_clock u2.mem\[63\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10345_ _04893_ u2.mem\[52\]\[3\] _04966_ _04970_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12007__D net25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10804__S _05253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13192__CLK clknet_leaf_276_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13064_ _00943_ clknet_leaf_47_clock u2.mem\[58\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10276_ _04930_ _00807_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12015_ net29 clknet_2_2__leaf_clock_a mem_address_trans\[5\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08231__I0 _03579_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07734__A2 _03013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12917_ _00796_ clknet_leaf_83_clock u2.mem\[49\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12848_ _00727_ clknet_leaf_151_clock u2.mem\[45\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_202_clock_I clknet_5_29_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12779_ _00658_ clknet_leaf_253_clock u2.mem\[41\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09839__I _04440_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08743__I _03962_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_159_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07359__I _02569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09798__I0 _04612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13535__CLK clknet_leaf_329_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07422__B2 u2.mem\[20\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09990_ _04752_ _00699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07973__A2 _02559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08941_ _04037_ u2.mem\[19\]\[10\] _04084_ _04087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11357__I0 _05593_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08222__I0 _03570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08872_ _03718_ _04046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07094__I _02572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07725__A2 _03080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07823_ u2.mem\[60\]\[12\] _03288_ _03289_ u2.mem\[62\]\[12\] _03290_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11545__S _05722_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07754_ u2.mem\[43\]\[11\] _03049_ _03050_ u2.mem\[20\]\[11\] _03222_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08918__I _04073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07822__I _02548_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06705_ u2.mem\[165\]\[1\] _02076_ _02079_ u2.mem\[163\]\[1\] _02092_ u2.mem\[177\]\[1\]
+ _02189_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_07685_ u2.mem\[5\]\[9\] _03153_ _03154_ u2.mem\[38\]\[9\] _03155_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11344__I _05516_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09424_ _04400_ _00485_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06636_ _02120_ _02121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08854__S _04033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06161__A1 u2.mem\[180\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06161__B2 u2.mem\[150\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09355_ _04353_ _00463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06567_ _01990_ _02032_ _02052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08306_ _03680_ _03681_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09286_ _04246_ u2.mem\[27\]\[0\] _04313_ _04314_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06498_ _01979_ _01924_ _01970_ _01980_ _01983_ _01464_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_165_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07661__A1 _03105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08237_ _03632_ _03633_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06464__A2 _01942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07269__I _02358_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09789__I0 _04599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09685__S _04554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06173__I _01679_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08168_ _03591_ _00038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07119_ _02597_ _02598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10624__S _05141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12902__CLK clknet_leaf_74_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08099_ mem_address_trans\[0\].data_sync _03543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10130_ _04817_ u2.mem\[46\]\[15\] _04835_ _04839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10061_ _04795_ u2.mem\[45\]\[5\] _04793_ _04796_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08213__I0 _03561_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_151_clock_I clknet_5_25_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10020__I0 _04696_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09961__I0 _04712_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10963_ _05335_ u2.mem\[135\]\[0\] _05356_ _05357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13408__CLK clknet_leaf_304_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12702_ _00581_ clknet_leaf_256_clock u2.mem\[36\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06688__C1 u2.mem\[193\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08764__S _03973_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10894_ _05311_ _01044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12633_ _00512_ clknet_leaf_103_clock u2.mem\[31\]\[14\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10087__I0 _04813_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08563__I _03835_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12564_ _00443_ clknet_leaf_95_clock u2.mem\[27\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_11_0_clock clknet_4_5_0_clock clknet_5_11_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__12432__CLK clknet_leaf_159_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11823__I1 u2.mem\[188\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11515_ _05671_ u2.mem\[169\]\[2\] _05700_ _05703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_76_clock_I clknet_5_8_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06455__A2 _01942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12495_ _00374_ clknet_leaf_163_clock u2.mem\[23\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07179__I _02525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09595__S _04506_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11446_ _05629_ u2.mem\[165\]\[2\] _05655_ _05658_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06207__A2 _01619_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12582__CLK clknet_leaf_100_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10534__S _05083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11377_ _05285_ _05606_ _05615_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_158_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09394__I _04160_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13116_ _00995_ clknet_leaf_261_clock u2.mem\[62\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10328_ _04913_ u2.mem\[51\]\[12\] _04959_ _04960_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11339__I0 _05591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07128__B _02434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08204__I0 _03552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13047_ _00926_ clknet_leaf_44_clock u2.mem\[57\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10259_ _04614_ _04920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08939__S _04084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07707__A2 _03120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10011__I0 _04687_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09952__I0 _04703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10711__A1 _03904_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06391__A1 u2.mem\[159\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07642__I _02504_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06391__B2 u2.mem\[149\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09704__I0 _04570_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13088__CLK clknet_leaf_245_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11511__I0 _05663_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07470_ u2.mem\[44\]\[6\] _02887_ _02888_ u2.mem\[42\]\[6\] _02943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08674__S _03915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_353_clock_I clknet_5_1_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07340__B1 _02661_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06421_ _01911_ _01922_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07891__A1 _03353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09140_ _04219_ _00382_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08473__I _03777_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06352_ u2.mem\[158\]\[4\] _01728_ _01729_ u2.mem\[151\]\[4\] _01732_ u2.mem\[168\]\[4\]
+ _01855_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_124_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07238__A4 _02714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09071_ _03581_ _03750_ _04179_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06283_ _01785_ _01786_ _01787_ _01788_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12925__CLK clknet_leaf_257_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07089__I _02363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08022_ mem_address_trans\[2\].data_sync mem_address_trans\[3\].data_sync _03483_
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_129_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06997__A3 _02446_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11578__I0 _05713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10444__S _05035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09973_ _04687_ u2.mem\[43\]\[2\] _04740_ _04743_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08924_ _04077_ _00308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10002__I0 _04716_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09943__I0 _04694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08855_ _04034_ _00282_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11750__I0 _05825_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12305__CLK clknet_leaf_164_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07806_ _02488_ _03273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08786_ _03989_ _03990_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08648__I _03656_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05998_ _01505_ row_col_select_trans.data_sync _01506_ _01507_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06382__B2 u2.mem\[183\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input13_I data_in_a[15] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_07737_ u2.mem\[40\]\[11\] _03018_ _03019_ u2.mem\[30\]\[11\] _03205_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09171__I1 u2.mem\[24\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12110__D _05992_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07668_ _03134_ _03135_ _03136_ _03137_ _03138_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_81_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12455__CLK clknet_leaf_127_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09407_ _04173_ _04389_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06619_ _02026_ _02011_ _02104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07882__A1 u2.mem\[14\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06685__A2 _02168_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07599_ _02581_ _03070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07882__B2 u2.mem\[12\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09338_ _04265_ u2.mem\[28\]\[6\] _04341_ _04344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07634__A1 u2.mem\[27\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06437__A2 _01915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09269_ _04274_ u2.mem\[26\]\[10\] _04300_ _04303_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11300_ _05567_ _05568_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_5_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12280_ _00159_ clknet_leaf_120_clock u2.mem\[9\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11231_ _05514_ u2.mem\[151\]\[4\] _05519_ _05525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08434__I0 _03710_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10241__I0 _04907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08985__I1 u2.mem\[20\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11162_ _05470_ u2.mem\[147\]\[4\] _05474_ _05480_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10113_ _04829_ _00745_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11093_ _05437_ _01117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08759__S _03968_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09934__I0 _04685_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10044_ _04783_ _04784_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_96_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11741__I0 _05833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11185__S _05492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13230__CLK clknet_leaf_279_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08362__A2 _03606_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06373__A1 _01848_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07570__B1 _03040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11995_ _00007_ clknet_leaf_319_clock u2.mem\[0\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08494__S _03800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10946_ _05343_ u2.mem\[134\]\[2\] _05337_ _05344_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07873__A1 u2.mem\[16\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06676__A2 _02142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10877_ _05299_ u2.mem\[130\]\[1\] _05297_ _05300_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12616_ _00495_ clknet_leaf_113_clock u2.mem\[30\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08293__I _03502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12547_ _00426_ clknet_leaf_103_clock u2.mem\[26\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12478_ _00357_ clknet_leaf_181_clock u2.mem\[22\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_304_clock clknet_5_16_0_clock clknet_leaf_304_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_67_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08425__I0 _03693_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11429_ _05648_ _01242_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10264__S _04923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08976__I1 u2.mem\[20\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11980__I0 _05222_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12328__CLK clknet_leaf_126_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06970_ u2.mem\[45\]\[0\] _02444_ _02448_ u2.mem\[34\]\[0\] _02449_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_319_clock clknet_5_18_0_clock clknet_leaf_319_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09925__I0 _04714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I col_select_a[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08640_ _03826_ u2.mem\[12\]\[12\] _03895_ _03896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06364__A1 u2.mem\[154\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12478__CLK clknet_leaf_181_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07372__I _02600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06364__B2 u2.mem\[162\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08571_ _03855_ _00177_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11823__S _05887_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07522_ u2.mem\[37\]\[7\] _02825_ _02826_ u2.mem\[59\]\[7\] _02994_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_165_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06116__A1 _01571_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07453_ _02905_ _02912_ _02919_ _02926_ _02927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__07864__A1 _03297_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06667__A2 _01999_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10439__S _05030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06404_ u2.mem\[146\]\[5\] _01691_ _01693_ u2.mem\[186\]\[5\] _01906_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_10_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06716__I _02137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07384_ _02613_ _02859_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09123_ _04145_ u2.mem\[23\]\[5\] _04208_ _04210_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06335_ _01836_ _01837_ _01838_ _01839_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08664__I0 _03912_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09054_ data_in_trans\[12\].data_sync _04166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07092__A2 _02565_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06266_ u2.mem\[171\]\[2\] _01611_ _01770_ u2.mem\[157\]\[2\] _01771_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_15_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13103__CLK clknet_leaf_312_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08005_ _01591_ _03464_ _03467_ _01678_ _03468_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__08416__I0 _03676_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10174__S _04865_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06197_ _01552_ _01615_ _01704_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07547__I _02405_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09963__S _04734_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07919__A2 _02503_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08967__I1 u2.mem\[20\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06451__I _01923_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11971__I0 _05213_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13253__CLK clknet_leaf_291_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09956_ _04707_ u2.mem\[42\]\[11\] _04729_ _04733_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08907_ _04041_ u2.mem\[18\]\[12\] _04066_ _04067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09887_ _04688_ _00660_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_24_clock_I clknet_5_2_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09392__I1 u2.mem\[29\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08838_ _04022_ _00277_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10701__I _05173_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06355__A1 u2.mem\[175\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06355__B2 u2.mem\[188\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07552__B1 _03022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08769_ _03977_ _00253_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10800_ _04416_ _05172_ _05252_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11780_ _05867_ _01374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07304__B1 _02758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10731_ _03683_ _05209_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06658__A2 _02077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11651__A2 _05769_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_249_clock_I clknet_5_22_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13450_ _01329_ clknet_leaf_343_clock u2.mem\[178\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10662_ _05166_ _00957_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11995__CLK clknet_leaf_319_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12401_ _00280_ clknet_leaf_161_clock u2.mem\[17\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08655__I0 _03900_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13381_ _01260_ clknet_leaf_305_clock u2.mem\[167\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10593_ _05126_ u2.mem\[57\]\[14\] _05122_ _05127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12332_ _00211_ clknet_leaf_206_clock u2.mem\[13\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10462__I0 _05020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07083__A2 _02559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06291__B1 _01715_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12263_ _00142_ clknet_leaf_55_clock u2.mem\[8\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08407__I0 _03657_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_301_clock_I clknet_5_16_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11167__A1 _04094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08958__I1 u2.mem\[20\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11214_ _05513_ _05514_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12194_ _00073_ clknet_leaf_238_clock u2.mem\[4\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11962__I0 _05913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_290_clock clknet_5_20_0_clock clknet_leaf_290_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__12015__D net29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11145_ _05469_ _01137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12620__CLK clknet_leaf_190_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11076_ _05342_ _05426_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09532__A1 _04013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10027_ _04703_ u2.mem\[44\]\[9\] _04772_ _04774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08288__I _03499_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06346__A1 u2.mem\[178\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07543__B1 _02867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06346__B2 u2.mem\[164\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12770__CLK clknet_leaf_155_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11978_ _05220_ u2.mem\[194\]\[11\] _05985_ _05987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06649__A2 _02033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10929_ _05331_ _01059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12000__CLK clknet_leaf_28_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08952__S _04089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13126__CLK clknet_leaf_23_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08646__I0 _03833_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10453__I0 _05011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06120_ _01621_ _01624_ _01626_ _01627_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_34_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_243_clock clknet_5_19_0_clock clknet_leaf_243_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_117_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12150__CLK clknet_leaf_73_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06051_ col_select_trans\[2\].data_sync _01558_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10205__I0 _04815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06271__I _01623_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11953__I0 _05903_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_258_clock clknet_5_23_0_clock clknet_leaf_258_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_114_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09810_ _04576_ u2.mem\[39\]\[3\] _04639_ _04643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10722__S _05196_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09741_ _04598_ _04599_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06953_ _02373_ _02432_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11705__I0 _05792_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_198_clock_I clknet_5_30_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09672_ _04476_ u2.mem\[36\]\[5\] _04549_ _04551_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06884_ _02362_ _02363_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08623_ _03886_ _00198_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06888__A2 _02338_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08554_ _03835_ _03846_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_39_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07505_ u2.mem\[16\]\[7\] _02798_ _02799_ u2.mem\[33\]\[7\] _02977_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07837__A1 u2.mem\[9\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08485_ _03798_ u2.mem\[9\]\[0\] _03800_ _03801_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_250_clock_I clknet_5_22_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07436_ u2.mem\[9\]\[5\] _02836_ _02837_ u2.mem\[25\]\[5\] _02910_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_11_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06446__I _01927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07367_ _02832_ _02835_ _02838_ _02841_ _02842_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08637__I0 _03824_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09106_ _04174_ u2.mem\[22\]\[14\] _04197_ _04200_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09757__I data_in_trans\[14\].data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10444__I0 _05001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06318_ u2.mem\[145\]\[3\] _01640_ _01732_ u2.mem\[168\]\[3\] _01822_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07298_ u2.mem\[5\]\[3\] _02687_ _02688_ u2.mem\[38\]\[3\] _02774_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09037_ data_in_trans\[8\].data_sync _04153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06249_ u2.mem\[166\]\[1\] _01753_ _01754_ u2.mem\[161\]\[1\] _01755_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12643__CLK clknet_leaf_94_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11944__I0 _05225_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06576__A1 _02058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07773__B1 _03089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09939_ _04723_ _00677_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07226__B _02359_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12950_ _00829_ clknet_leaf_30_clock u2.mem\[51\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06328__A1 u2.mem\[152\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07525__B1 _02907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11901_ u2.mem\[192\]\[10\] _03523_ _05942_ _05943_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12881_ _00760_ clknet_leaf_143_clock u2.mem\[47\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07540__A3 _03006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11832_ _05899_ _01394_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08836__I _03671_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12023__CLK clknet_2_1__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13149__CLK clknet_leaf_264_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08876__I0 _04048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11763_ _05856_ _05857_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_26_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13502_ _01381_ clknet_leaf_331_clock u2.mem\[187\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10714_ _05197_ _00978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11694_ _05814_ _01341_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13433_ _01312_ clknet_leaf_338_clock u2.mem\[175\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08628__I0 _03815_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12173__CLK clknet_leaf_210_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13299__CLK clknet_leaf_363_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10645_ _05151_ _05157_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_35_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10435__I0 _04987_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13364_ _01243_ clknet_leaf_358_clock u2.mem\[164\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10576_ _03696_ _05115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12315_ _00194_ clknet_leaf_222_clock u2.mem\[12\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13295_ _01174_ clknet_leaf_2_clock u2.mem\[152\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12246_ _00125_ clknet_leaf_73_clock u2.mem\[7\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08005__A1 _01591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08005__B2 _01678_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11935__I0 _05216_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11638__S _05779_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08800__I0 _03919_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12177_ _00056_ clknet_leaf_218_clock u2.mem\[3\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07764__B1 _03070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09108__S _04197_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11128_ _05430_ u2.mem\[145\]\[4\] _05452_ _05458_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11059_ _05415_ _01105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07516__B1 _02894_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06319__B2 u2.mem\[188\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11373__S _05607_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07650__I _02520_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07819__A1 _03257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08867__I0 _04041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08270_ _03652_ _00079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07295__A2 _02601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07221_ u2.mem\[27\]\[2\] _02428_ _02436_ u2.mem\[35\]\[2\] _02698_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_182_clock clknet_5_27_0_clock clknet_leaf_182_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08619__I0 _03806_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11900__I _05927_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07152_ _02615_ _02620_ _02625_ _02630_ _02631_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_34_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09292__I0 _04258_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12666__CLK clknet_leaf_56_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06103_ _01607_ _01609_ _01610_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07083_ u2.mem\[61\]\[0\] _02559_ _02561_ u2.mem\[63\]\[0\] _02562_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_197_clock clknet_5_30_0_clock clknet_leaf_197_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_12_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06034_ inverter_select_trans.data_sync _01542_ _01543_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09044__I0 _04158_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11926__I0 _05915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10729__I1 u2.mem\[61\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07825__I _02541_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_120_clock clknet_5_15_0_clock clknet_leaf_120_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07985_ u2.mem\[52\]\[15\] _03313_ _03314_ u2.mem\[21\]\[15\] _03449_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09347__I1 u2.mem\[28\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09724_ _04585_ _04586_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06936_ _02414_ _02415_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07046__B _02411_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08857__S _04033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11154__I1 u2.mem\[147\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09655_ _04540_ _00576_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06867_ _02338_ _02345_ _02346_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08606_ _03875_ _00192_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_135_clock clknet_5_13_0_clock clknet_leaf_135_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09586_ _04463_ u2.mem\[34\]\[0\] _04501_ _04502_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07560__I _02474_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06730__A1 u2.mem\[180\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06798_ u2.mem\[167\]\[4\] _02059_ _02061_ u2.mem\[183\]\[4\] _02279_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08537_ _03798_ u2.mem\[10\]\[0\] _03836_ _03837_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12196__CLK clknet_leaf_71_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11606__A2 _05729_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11082__I _05348_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13441__CLK clknet_leaf_348_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08592__S _03867_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08468_ _03790_ _00139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07286__A2 _02554_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07419_ _02530_ _02893_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08399_ _03747_ _00113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11810__I _05768_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08391__I _03727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10430_ _03721_ _05027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06904__I _02351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11090__I0 _05420_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10361_ _04909_ u2.mem\[52\]\[10\] _04976_ _04979_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06797__A1 u2.mem\[164\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12100_ _01498_ clknet_leaf_149_clock u2.active_mem\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06797__B2 u2.mem\[178\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09035__I0 _04151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13080_ _00959_ clknet_leaf_43_clock u2.mem\[59\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10292_ _04939_ _00814_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06261__A3 _01758_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11917__I0 _05907_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12031_ net40 clknet_2_3__leaf_clock_a row_select_trans\[3\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09586__I1 u2.mem\[34\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06549__A1 _02031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07746__B1 _03112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12933_ _00812_ clknet_leaf_67_clock u2.mem\[50\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07513__A3 _02983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12864_ _00743_ clknet_leaf_148_clock u2.mem\[46\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06721__A1 _01727_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06721__B2 _02204_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11815_ _05868_ u2.mem\[188\]\[1\] _05888_ _05890_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12795_ _00674_ clknet_leaf_220_clock u2.mem\[42\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11921__S _05950_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07277__A2 _02654_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11746_ _05846_ _01361_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_146_clock_I clknet_5_24_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11677_ _05804_ _01334_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09397__I _04163_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10628_ _05147_ _00942_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13416_ _01295_ clknet_leaf_341_clock u2.mem\[172\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09274__I0 _04278_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10336__I _04862_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13347_ _01226_ clknet_leaf_17_clock u2.mem\[161\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10559_ _05000_ _05103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13278_ _01157_ clknet_leaf_9_clock u2.mem\[149\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12229_ _00108_ clknet_leaf_69_clock u2.mem\[6\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12069__CLK clknet_2_0__leaf_clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07645__I _02510_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13314__CLK clknet_leaf_349_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09329__I1 u2.mem\[28\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07770_ u2.mem\[18\]\[11\] _03083_ _03084_ u2.mem\[19\]\[11\] _03238_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08677__S _03915_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_52_clock clknet_5_12_0_clock clknet_leaf_52_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06721_ _01727_ _01995_ _02171_ _02204_ _01475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09440_ _04409_ _00492_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13464__CLK clknet_leaf_344_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06652_ _02006_ _02002_ _02137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10895__I0 _05299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07380__I _02616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09371_ _04135_ _04364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06583_ _02067_ _02068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_67_clock clknet_5_9_0_clock clknet_leaf_67_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_40_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11831__S _05896_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08322_ _03659_ _03694_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_75_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07268__A2 _02475_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08253_ _03559_ u2.mem\[4\]\[6\] _03640_ _03643_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07204_ u2.mem\[23\]\[1\] _02680_ _02681_ u2.mem\[22\]\[1\] _02682_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09265__I0 _04269_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08184_ _03584_ _03600_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_118_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07135_ _02613_ _02614_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06779__A1 u2.mem\[180\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06779__B2 u2.mem\[172\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07066_ _02544_ _02537_ _02538_ _02519_ _02545_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_134_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_348_clock_I clknet_5_4_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06017_ u2.driver_mem\[4\] _01517_ _01525_ _01520_ _01526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_160_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07728__B1 _03154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11524__A1 _04287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07555__I _02460_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09971__S _04740_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06400__B1 _01672_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07968_ u2.mem\[14\]\[15\] _02526_ _02528_ u2.mem\[12\]\[15\] _03432_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10910__S _05319_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06919_ _02363_ _02398_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09707_ _04572_ _04573_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07899_ u2.mem\[52\]\[13\] _03313_ _03314_ u2.mem\[21\]\[13\] _03365_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10886__I0 _05305_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09638_ _04480_ u2.mem\[35\]\[7\] _04527_ _04531_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09569_ _04489_ u2.mem\[33\]\[11\] _04483_ _04490_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11741__S _05840_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11600_ _05676_ _05756_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12580_ _00459_ clknet_leaf_98_clock u2.mem\[28\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07259__A2 _02725_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11531_ _05670_ _05713_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10357__S _04976_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12981__CLK clknet_leaf_31_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11462_ _05668_ u2.mem\[166\]\[1\] _05665_ _05669_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09256__I0 _04260_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09010__I _04131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13201_ _01080_ clknet_leaf_278_clock u2.mem\[137\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10413_ _05015_ _00859_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11393_ _05624_ _05625_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07967__B1 _02523_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13132_ _01011_ clknet_leaf_267_clock u2.mem\[63\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10344_ _04969_ _00836_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13337__CLK clknet_leaf_9_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07431__A2 _02902_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13063_ _00942_ clknet_leaf_48_clock u2.mem\[58\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10275_ _04898_ u2.mem\[50\]\[5\] _04928_ _04930_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07719__B1 _03067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12014_ mem_address_trans\[4\].A clknet_leaf_289_clock mem_address_trans\[4\].data_sync
+ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12361__CLK clknet_leaf_133_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10820__S _05263_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_72_clock_I clknet_5_8_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10877__I0 _05299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12916_ _00795_ clknet_leaf_60_clock u2.mem\[49\]\[9\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07498__A2 _02866_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12847_ _00726_ clknet_leaf_151_clock u2.mem\[45\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10629__I0 _05124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_12778_ _00657_ clknet_leaf_130_clock u2.mem\[40\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_297_clock_I clknet_5_17_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11729_ _05836_ _01354_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09247__I0 _04246_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08960__S _04097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10066__I _04588_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11098__S _05434_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08940_ _04086_ _00315_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12704__CLK clknet_leaf_238_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07375__I _02605_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09791__S _04628_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11357__I1 u2.mem\[159\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_08871_ _04045_ _00287_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07822_ _02548_ _03289_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12854__CLK clknet_leaf_80_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07753_ u2.mem\[49\]\[11\] _03126_ _03127_ u2.mem\[46\]\[11\] _03221_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08200__S _03609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06704_ u2.mem\[188\]\[1\] _02185_ _02186_ u2.mem\[187\]\[1\] _02187_ u2.mem\[192\]\[1\]
+ _02188_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__10868__I0 _05207_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07684_ _02628_ _03154_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09423_ _04364_ u2.mem\[30\]\[3\] _04396_ _04400_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06635_ _02119_ _02000_ _02120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09354_ _04281_ u2.mem\[28\]\[13\] _04351_ _04353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06566_ _02050_ _02051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08305_ _03679_ _03680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09285_ _04312_ _04313_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06497_ u2.mem\[193\]\[15\] _01917_ _01982_ _01911_ _01983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_20_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08236_ _03631_ mem_address_trans\[3\].data_sync _03632_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09238__I0 _04283_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08870__S _04042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12234__CLK clknet_leaf_52_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06454__I _01913_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07661__A2 _03110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11045__I0 _05386_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08167_ _03554_ u2.mem\[2\]\[4\] _03590_ _03591_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09789__I1 u2.mem\[38\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07118_ _02418_ _02420_ _02507_ _02426_ _02597_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_88_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08098_ _03541_ _03542_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12384__CLK clknet_leaf_221_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06621__B1 _02105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07049_ _02527_ _02528_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10060_ _04582_ _04795_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09206__S _04261_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10962_ _05355_ _05356_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_28_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09005__I _04127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12701_ _00580_ clknet_leaf_257_clock u2.mem\[36\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06688__C2 _02089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_10893_ _05294_ u2.mem\[131\]\[0\] _05310_ _05311_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12632_ _00511_ clknet_leaf_104_clock u2.mem\[31\]\[13\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12563_ _00442_ clknet_leaf_94_clock u2.mem\[27\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11514_ _05702_ _01273_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_19_clock_I clknet_5_2_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12494_ _00373_ clknet_leaf_181_clock u2.mem\[23\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07652__A2 _03120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11036__I0 _05392_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12018__D mem_address_trans\[6\].A vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11445_ _05657_ _01249_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12727__CLK clknet_leaf_43_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11376_ _05614_ _01223_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10327_ _04943_ _04959_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_13115_ _00994_ clknet_5_22_0_clock u2.mem\[62\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07195__I _02572_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11339__I1 u2.mem\[158\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13046_ _00925_ clknet_leaf_25_clock u2.mem\[57\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_10258_ _04919_ _00800_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12877__CLK clknet_leaf_214_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07128__C _02483_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11646__S _05778_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10189_ _04799_ u2.mem\[48\]\[7\] _04870_ _04874_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09116__S _04203_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12107__CLK clknet_leaf_135_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06391__A2 _01603_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09704__I1 u2.mem\[37\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11511__I1 u2.mem\[169\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11381__S _05616_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06420_ u2.mem\[193\]\[0\] _01917_ _01919_ u2.mem\[192\]\[0\] _01920_ _01921_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_22_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12257__CLK clknet_leaf_228_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13502__CLK clknet_leaf_331_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06351_ u2.mem\[145\]\[4\] _01639_ _01643_ u2.mem\[163\]\[4\] u2.mem\[165\]\[4\]
+ _01645_ _01854_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_72_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09070_ _04178_ _00353_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08690__S _03924_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06282_ u2.mem\[159\]\[2\] _01604_ _01595_ u2.mem\[149\]\[2\] _01787_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07643__A2 _03111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08021_ mem_address_trans\[0\].data_sync _03482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_159_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06851__B1 _02147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06997__A4 _02463_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09585__I _04500_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09972_ _04742_ _00691_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08923_ _04019_ u2.mem\[19\]\[2\] _04074_ _04077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07159__B2 u2.mem\[30\]\[1\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08854_ _04032_ u2.mem\[17\]\[8\] _04033_ _04034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06906__A1 _02364_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07833__I _02569_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11750__I1 u2.mem\[184\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07805_ _02485_ _03272_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_08785_ _03983_ _03988_ _03989_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_22_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05997_ u2.select_mem_row\[0\] row_col_select_trans.data_sync _01506_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13032__CLK clknet_leaf_328_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07736_ u2.mem\[32\]\[11\] _03015_ _03016_ u2.mem\[2\]\[11\] _03204_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07667_ u2.mem\[57\]\[9\] _03061_ _03062_ u2.mem\[41\]\[9\] _03137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09406_ _04388_ _00479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06618_ _02053_ _02012_ _02103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07598_ _02579_ _03069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07882__A2 _02526_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13182__CLK clknet_leaf_271_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09337_ _04343_ _00455_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06549_ _02031_ _02033_ _02034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_20_clock_I clknet_5_2_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09268_ _04302_ _00427_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07634__A2 _03021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08219_ _03621_ _00059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09199_ _04256_ u2.mem\[25\]\[2\] _04252_ _04257_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09495__I _04442_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11230_ _05524_ _01167_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08434__I1 u2.mem\[7\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11161_ _05479_ _01143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10434__I _05029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10112_ _04799_ u2.mem\[46\]\[7\] _04825_ _04829_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06070__A1 _01552_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11092_ _05424_ u2.mem\[143\]\[1\] _05435_ _05437_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_245_clock_I clknet_5_22_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08198__I0 _03539_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10043_ _03904_ _04760_ _04783_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_49_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08839__I _03675_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07743__I _02357_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11741__I1 u2.mem\[183\]\[3\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06373__A2 _01853_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08775__S _03978_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11994_ _00006_ clknet_leaf_320_clock u2.mem\[0\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10945_ _05342_ _05343_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06125__A2 _01609_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10876_ _04991_ _05299_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12615_ _00494_ clknet_leaf_113_clock u2.mem\[30\]\[12\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08122__I0 _03559_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12546_ _00425_ clknet_leaf_168_clock u2.mem\[26\]\[7\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07625__A2 _03094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12477_ _00356_ clknet_leaf_181_clock u2.mem\[22\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11428_ _05623_ u2.mem\[164\]\[0\] _05647_ _05648_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08425__I1 u2.mem\[7\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11359_ _05595_ u2.mem\[159\]\[5\] _05597_ _05604_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08189__I0 _03577_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13055__CLK clknet_leaf_240_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_13029_ _00908_ clknet_leaf_31_clock u2.mem\[56\]\[10\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07653__I _02525_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06364__A2 _01699_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08570_ _03833_ u2.mem\[10\]\[15\] _03851_ _03855_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07521_ u2.mem\[60\]\[7\] _02822_ _02823_ u2.mem\[62\]\[7\] _02993_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06116__A2 _01617_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07452_ _02922_ _02923_ _02924_ _02925_ _02926_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08484__I _03799_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07864__A2 _03308_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06403_ u2.mem\[191\]\[5\] _01681_ _01683_ u2.mem\[179\]\[5\] _01905_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11248__I0 _05517_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_07383_ _02611_ _02858_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09122_ _04209_ _00374_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06334_ u2.mem\[146\]\[3\] _01692_ _01694_ u2.mem\[186\]\[3\] _01838_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07616__A2 _02920_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_194_clock_I clknet_5_31_0_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_09053_ _04165_ _00349_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06265_ _01614_ _01770_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10455__S _05040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08004_ _03465_ _03466_ _03467_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07828__I _02555_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09613__I0 _04491_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_06196_ _01702_ _01703_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11971__I1 u2.mem\[194\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09955_ _04732_ _00684_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08906_ _04050_ _04066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_131_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09886_ _04687_ u2.mem\[41\]\[2\] _04683_ _04688_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07563__I _02479_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08837_ _04021_ u2.mem\[17\]\[3\] _04015_ _04022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07552__A1 u2.mem\[27\]\[8\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11085__I _05351_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06355__A2 _01601_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08768_ _03930_ u2.mem\[15\]\[11\] _03973_ _03977_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07719_ u2.mem\[29\]\[10\] _03066_ _03067_ u2.mem\[11\]\[10\] _03188_ vccd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07304__A1 _01808_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06107__A2 _01612_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08699_ _03718_ _03937_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10730_ _05208_ _00983_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06907__I _02385_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10661_ _05119_ u2.mem\[59\]\[11\] _05162_ _05166_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12400_ _00279_ clknet_leaf_156_clock u2.mem\[17\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13380_ _01259_ clknet_leaf_352_clock u2.mem\[166\]\[5\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10592_ _03717_ _05126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12331_ _00210_ clknet_leaf_207_clock u2.mem\[13\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06291__A1 u2.mem\[152\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_12262_ _00141_ clknet_leaf_69_clock u2.mem\[8\]\[11\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09604__I0 _04482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06291__B2 u2.mem\[148\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11167__A2 _05482_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13078__CLK clknet_leaf_25_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_11213_ _03506_ _05513_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12193_ _00072_ clknet_leaf_228_clock u2.mem\[4\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11144_ _05468_ u2.mem\[146\]\[3\] _05462_ _05469_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11962__I1 u2.mem\[194\]\[4\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07240__B1 _02549_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11075_ _05425_ _01111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10026_ _04773_ _00714_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09532__A2 _04441_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11924__S _05955_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12031__D net40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12915__CLK clknet_leaf_147_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06089__I _01587_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11478__I0 _05680_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_11977_ _05986_ _01452_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10928_ _05303_ u2.mem\[133\]\[3\] _05327_ _05331_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_0_clock_a_I clock_a vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10859_ _05288_ _01032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08646__I1 u2.mem\[12\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_13578_ _01457_ clknet_leaf_37_clock u2.mem\[194\]\[15\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12529_ _00408_ clknet_leaf_166_clock u2.mem\[25\]\[6\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06050_ _01556_ _01557_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06282__A1 u2.mem\[159\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06282__B2 u2.mem\[149\]\[2\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06034__A1 inverter_select_trans.data_sync vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12445__CLK clknet_leaf_198_clock vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11953__I1 u2.mem\[194\]\[0\] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09740_ data_in_trans\[10\].data_sync _04598_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06952_ _02430_ _02431_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_113_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
.ends

